
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER
-- DATE: Mon May 14 10:21:16 2018

	signal mem : ram_t := (  -- TODO: Promeniti velicinu mem. Choice 8192 is out of range 0 to 8191 for the index subtype.
	
	--			***** COLOR PALLETE *****

		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00000700", -- R: 0 G: 7 B: 0
		2 =>	x"0000077D", -- R: 125 G: 7 B: 0
		3 =>	x"003C0000", -- R: 0 G: 0 B: 60
		4 =>	x"00D8AC4A", -- R: 74 G: 172 B: 216
		5 =>	x"00006092", -- R: 146 G: 96 B: 0
		6 =>	x"00460000", -- R: 0 G: 0 B: 70
		7 =>	x"000C0000", -- R: 0 G: 0 B: 12
		8 =>	x"000C7D3C", -- R: 60 G: 125 B: 12
		9 =>	x"00000070", -- R: 112 G: 0 B: 0
		10 =>	x"00AC4A00", -- R: 0 G: 74 B: 172
		11 =>	x"0068C04A", -- R: 74 G: 192 B: 104
		12 =>	x"006D005C", -- R: 92 G: 0 B: 109
		13 =>	x"00006200", -- R: 0 G: 98 B: 0
		14 =>	x"0069006E", -- R: 110 G: 0 B: 105
		15 =>	x"00005C00", -- R: 0 G: 92 B: 0
		16 =>	x"00310036", -- R: 54 G: 0 B: 49
		17 =>	x"00007800", -- R: 0 G: 120 B: 0
		18 =>	x"00620061", -- R: 97 G: 0 B: 98
		19 =>	x"00006E00", -- R: 0 G: 110 B: 0
		20 =>	x"0067002E", -- R: 46 G: 0 B: 103
		21 =>	x"006D0070", -- R: 112 G: 0 B: 109
		22 =>	x"005C0062", -- R: 98 G: 0 B: 92
		23 =>	x"00006300", -- R: 0 G: 99 B: 0
		24 =>	x"005F006D", -- R: 109 G: 0 B: 95
		25 =>	x"00006500", -- R: 0 G: 101 B: 0
		26 =>	x"006D005F", -- R: 95 G: 0 B: 109
		27 =>	x"00007000", -- R: 0 G: 112 B: 0
		28 =>	x"00610063", -- R: 99 G: 0 B: 97
		29 =>	x"00006B00", -- R: 0 G: 107 B: 0
		30 =>	x"00650072", -- R: 114 G: 0 B: 101
		31 =>	x"00007400", -- R: 0 G: 116 B: 0
		32 =>	x"0074006C", -- R: 108 G: 0 B: 116
		33 =>	x"00310035", -- R: 53 G: 0 B: 49
		34 =>	x"00310034", -- R: 52 G: 0 B: 49
		35 =>	x"00002D00", -- R: 0 G: 45 B: 0
		36 =>	x"0035002D", -- R: 45 G: 0 B: 53
		37 =>	x"00003200", -- R: 0 G: 50 B: 0
		38 =>	x"00300031", -- R: 49 G: 0 B: 48
		39 =>	x"00003800", -- R: 0 G: 56 B: 0
		40 =>	x"005C006E", -- R: 110 G: 0 B: 92
		41 =>	x"0077005F", -- R: 95 G: 0 B: 119
		42 =>	x"00007200", -- R: 0 G: 114 B: 0
		43 =>	x"0061006C", -- R: 108 G: 0 B: 97
		44 =>	x"00006C00", -- R: 0 G: 108 B: 0
		45 =>	x"0079005F", -- R: 95 G: 0 B: 121
		46 =>	x"0048104B", -- R: 75 G: 16 B: 72
		47 =>	x"0000D8AC", -- R: 172 G: 216 B: 0
		48 =>	x"004A0044", -- R: 68 G: 0 B: 74
		49 =>	x"00003A00", -- R: 0 G: 58 B: 0
		50 =>	x"005C006D", -- R: 109 G: 0 B: 92
		51 =>	x"00006100", -- R: 0 G: 97 B: 0
		52 =>	x"00740065", -- R: 101 G: 0 B: 116
		53 =>	x"0069006A", -- R: 106 G: 0 B: 105
		54 =>	x"005C0052", -- R: 82 G: 0 B: 92
		55 =>	x"00004100", -- R: 0 G: 65 B: 0
		56 =>	x"00320031", -- R: 49 G: 0 B: 50
		57 =>	x"002D0032", -- R: 50 G: 0 B: 45
		58 =>	x"00003000", -- R: 0 G: 48 B: 0
		59 =>	x"00DDDDDD", -- R: 221 G: 221 B: 221
		60 =>	x"00DDDD5C", -- R: 92 G: 221 B: 221
		61 =>	x"00004C00", -- R: 0 G: 76 B: 0
		62 =>	x"00004C24", -- R: 36 G: 76 B: 0
		63 =>	x"003FFE00", -- R: 0 G: 254 B: 63
		64 =>	x"00007CFE", -- R: 254 G: 124 B: 0
		65 =>	x"00000060", -- R: 96 G: 0 B: 0
		66 =>	x"00760000", -- R: 0 G: 0 B: 118
		67 =>	x"00002000", -- R: 0 G: 32 B: 0
		68 =>	x"0000FDFD", -- R: 253 G: 253 B: 0
		69 =>	x"00FDFDDD", -- R: 221 G: 253 B: 253
		70 =>	x"006CDDBF", -- R: 191 G: 221 B: 108
		71 =>	x"0045363C", -- R: 60 G: 54 B: 69
		72 =>	x"00000048", -- R: 72 G: 0 B: 0
		73 =>	x"00104B00", -- R: 0 G: 75 B: 16
		74 =>	x"0000DDDD", -- R: 221 G: 221 B: 0
		75 =>	x"00008000", -- R: 0 G: 128 B: 0
		76 =>	x"0000C0C0", -- R: 192 G: 192 B: 0
		77 =>	x"00000071", -- R: 113 G: 0 B: 0
		78 =>	x"00E00000", -- R: 0 G: 0 B: 224
		79 =>	x"007BF000", -- R: 0 G: 240 B: 123
		80 =>	x"0000156C", -- R: 108 G: 21 B: 0
		81 =>	x"00000015", -- R: 21 G: 0 B: 0
		82 =>	x"006A0000", -- R: 0 G: 0 B: 106
		83 =>	x"00156A00", -- R: 0 G: 106 B: 21
		84 =>	x"00003148", -- R: 72 G: 49 B: 0
		85 =>	x"002A0000", -- R: 0 G: 0 B: 42
		86 =>	x"00556800", -- R: 0 G: 104 B: 85
		87 =>	x"00005568", -- R: 104 G: 85 B: 0
		88 =>	x"0000003B", -- R: 59 G: 0 B: 0
		89 =>	x"006C0000", -- R: 0 G: 0 B: 108
		90 =>	x"00FF0000", -- R: 0 G: 0 B: 255
		91 =>	x"00FFFF00", -- R: 0 G: 255 B: 255
		92 =>	x"0000FFFF", -- R: 255 G: 255 B: 0
		93 =>	x"000000FF", -- R: 255 G: 0 B: 0
		94 =>	x"0000FF00", -- R: 0 G: 255 B: 0
		95 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		96 =>	x"00FF00FF", -- R: 255 G: 0 B: 255
		97 =>	x"004600D8", -- R: 216 G: 0 B: 70
		98 =>	x"00609246", -- R: 70 G: 146 B: 96
		99 =>	x"00000400", -- R: 0 G: 4 B: 0
		100 =>	x"0000047D", -- R: 125 G: 4 B: 0
		101 =>	x"006D0061", -- R: 97 G: 0 B: 109
		102 =>	x"005F0065", -- R: 101 G: 0 B: 95
		103 =>	x"0065006D", -- R: 109 G: 0 B: 101
		104 =>	x"006E0074", -- R: 116 G: 0 B: 110
		105 =>	x"00005F00", -- R: 0 G: 95 B: 0
		106 =>	x"00300030", -- R: 48 G: 0 B: 48
		107 =>	x"00002E00", -- R: 0 G: 46 B: 0
		108 =>	x"0062006D", -- R: 109 G: 0 B: 98
		109 =>	x"00DD3A00", -- R: 0 G: 58 B: 221
		110 =>	x"00004900", -- R: 0 G: 73 B: 0
		111 =>	x"00004927", -- R: 39 G: 73 B: 0
		112 =>	x"0050204B", -- R: 75 G: 32 B: 80
		113 =>	x"004A00DD", -- R: 221 G: 0 B: 74
		114 =>	x"00112000", -- R: 0 G: 32 B: 17
		115 =>	x"00220022", -- R: 34 G: 0 B: 34
		116 =>	x"00001111", -- R: 17 G: 17 B: 0
		117 =>	x"00302002", -- R: 2 G: 32 B: 48
		118 =>	x"00560011", -- R: 17 G: 0 B: 86
		119 =>	x"00111111", -- R: 17 G: 17 B: 17
		120 =>	x"00200202", -- R: 2 G: 2 B: 32
		121 =>	x"00031111", -- R: 17 G: 17 B: 3
		122 =>	x"00313311", -- R: 17 G: 51 B: 49
		123 =>	x"001111FD", -- R: 253 G: 17 B: 17
		124 =>	x"00FDFDFD", -- R: 253 G: 253 B: 253
		125 =>	x"00DD64DD", -- R: 221 G: 100 B: 221
		126 =>	x"00BF4D2E", -- R: 46 G: 77 B: 191
		127 =>	x"00300005", -- R: 5 G: 0 B: 48
		128 =>	x"00020020", -- R: 32 G: 0 B: 2
		129 =>	x"00202330", -- R: 48 G: 35 B: 32
		130 =>	x"00050000", -- R: 0 G: 0 B: 5
		131 =>	x"00033522", -- R: 34 G: 53 B: 3
		132 =>	x"00022322", -- R: 34 G: 35 B: 2
		133 =>	x"00024033", -- R: 51 G: 64 B: 2
		134 =>	x"00300000", -- R: 0 G: 0 B: 48
		135 =>	x"00020004", -- R: 4 G: 0 B: 2
		136 =>	x"00400332", -- R: 50 G: 3 B: 64
		137 =>	x"00200422", -- R: 34 G: 4 B: 32
		138 =>	x"00042000", -- R: 0 G: 32 B: 4
		139 =>	x"00031300", -- R: 0 G: 19 B: 3
		140 =>	x"00002204", -- R: 4 G: 34 B: 0
		141 =>	x"00222331", -- R: 49 G: 35 B: 34
		142 =>	x"00333311", -- R: 17 G: 51 B: 51
		143 =>	x"00113055", -- R: 85 G: 48 B: 17
		144 =>	x"00043111", -- R: 17 G: 49 B: 4
		145 =>	x"00111135", -- R: 53 G: 17 B: 17
		146 =>	x"00025022", -- R: 34 G: 80 B: 2
		147 =>	x"00002311", -- R: 17 G: 35 B: 0
		148 =>	x"00112002", -- R: 2 G: 32 B: 17
		149 =>	x"00002220", -- R: 32 G: 34 B: 0
		150 =>	x"00003110", -- R: 16 G: 49 B: 0
		151 =>	x"00022220", -- R: 32 G: 34 B: 2
		152 =>	x"00022022", -- R: 34 G: 32 B: 2
		153 =>	x"00313200", -- R: 0 G: 50 B: 49
		154 =>	x"00002042", -- R: 66 G: 32 B: 0
		155 =>	x"00002323", -- R: 35 G: 35 B: 0
		156 =>	x"009800FF", -- R: 255 G: 0 B: 152
		157 =>	x"00FF9800", -- R: 0 G: 152 B: 255
		158 =>	x"00FFFF98", -- R: 152 G: 255 B: 255
		159 =>	x"00A4FF98", -- R: 152 G: 255 B: 164
		160 =>	x"009800A4", -- R: 164 G: 0 B: 152
		161 =>	x"0000FF98", -- R: 152 G: 255 B: 0
		162 =>	x"0000A4FF", -- R: 255 G: 164 B: 0
		163 =>	x"00980000", -- R: 0 G: 0 B: 152
		164 =>	x"00A4FF99", -- R: 153 G: 255 B: 164
		165 =>	x"00980094", -- R: 148 G: 0 B: 152
		166 =>	x"00FF8621", -- R: 33 G: 134 B: 255
		167 =>	x"0036FF98", -- R: 152 G: 255 B: 54
		168 =>	x"000124FF", -- R: 255 G: 36 B: 1
		169 =>	x"00980095", -- R: 149 G: 0 B: 152
		170 =>	x"00A5FF98", -- R: 152 G: 255 B: 165
		171 =>	x"005480D7", -- R: 215 G: 128 B: 84
		172 =>	x"0038FF99", -- R: 153 G: 255 B: 56
		173 =>	x"009800DF", -- R: 223 G: 0 B: 152
		174 =>	x"0000DFFF", -- R: 255 G: 223 B: 0
		175 =>	x"0094FF99", -- R: 153 G: 255 B: 148
		176 =>	x"000095FF", -- R: 255 G: 149 B: 0
		177 =>	x"00980124", -- R: 36 G: 1 B: 152
		178 =>	x"00FF9900", -- R: 0 G: 153 B: 255
		179 =>	x"0000FF86", -- R: 134 G: 255 B: 0
		180 =>	x"002138FF", -- R: 255 G: 56 B: 33
		181 =>	x"0036FF99", -- R: 153 G: 255 B: 54
		182 =>	x"0000A7FF", -- R: 255 G: 167 B: 0
		183 =>	x"0098016B", -- R: 107 G: 1 B: 152
		184 =>	x"0038FF98", -- R: 152 G: 255 B: 56
		185 =>	x"00016BFF", -- R: 255 G: 107 B: 1
		186 =>	x"009800A7", -- R: 167 G: 0 B: 152
		187 =>	x"00320035", -- R: 53 G: 0 B: 50
		188 =>	x"0072006F", -- R: 111 G: 0 B: 114
		189 =>	x"006B002E", -- R: 46 G: 0 B: 107
		190 =>	x"00DD4C00", -- R: 0 G: 76 B: 221
		191 =>	x"00102000", -- R: 0 G: 32 B: 16
		192 =>	x"00000820", -- R: 32 G: 8 B: 0
		193 =>	x"00000007", -- R: 7 G: 0 B: 0
		194 =>	x"00C00000", -- R: 0 G: 0 B: 192
		195 =>	x"00000050", -- R: 80 G: 0 B: 0
		196 =>	x"00204B00", -- R: 0 G: 75 B: 32
		197 =>	x"001EC000", -- R: 0 G: 192 B: 30
		198 =>	x"00002020", -- R: 32 G: 32 B: 0
		199 =>	x"00000061", -- R: 97 G: 0 B: 0
		200 =>	x"00100000", -- R: 0 G: 0 B: 16
		201 =>	x"0081B000", -- R: 0 G: 176 B: 129
		202 =>	x"0000889E", -- R: 158 G: 136 B: 0
		203 =>	x"00000049", -- R: 73 G: 0 B: 0
		204 =>	x"00020000", -- R: 0 G: 0 B: 2
		205 =>	x"00CB0900", -- R: 0 G: 9 B: 203
		206 =>	x"0000890B", -- R: 11 G: 137 B: 0
		207 =>	x"000000BD", -- R: 189 G: 0 B: 0
		208 =>	x"00110000", -- R: 0 G: 0 B: 17
		209 =>	x"00610300", -- R: 0 G: 3 B: 97
		210 =>	x"0000271E", -- R: 30 G: 39 B: 0
		211 =>	x"00000030", -- R: 48 G: 0 B: 0
		212 =>	x"00600000", -- R: 0 G: 0 B: 96
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
		255 =>	x"00000000", -- Unused

--			***** 16x16 IMAGES *****

		256 =>	x"00000000", -- IMG_16x16_bang
		257 =>	x"00010203",
		258 =>	x"04050600",
		259 =>	x"00000000",
		260 =>	x"00000000",
		261 =>	x"00000000",
		262 =>	x"0708090A",
		263 =>	x"0B000000",
		264 =>	x"00000000",
		265 =>	x"00000000",
		266 =>	x"00000000",
		267 =>	x"00000000",
		268 =>	x"00000000",
		269 =>	x"00000000",
		270 =>	x"00000000",
		271 =>	x"00000000",
		272 =>	x"00000000",
		273 =>	x"00000000",
		274 =>	x"00000000",
		275 =>	x"00000000",
		276 =>	x"00000000",
		277 =>	x"00000000",
		278 =>	x"00000000",
		279 =>	x"00000000",
		280 =>	x"00000000",
		281 =>	x"00000000",
		282 =>	x"00000000",
		283 =>	x"00000000",
		284 =>	x"00000000",
		285 =>	x"00000000",
		286 =>	x"00000000",
		287 =>	x"00000000",
		288 =>	x"0C0D0E0F",
		289 =>	x"1011100F",
		290 =>	x"1213140D",
		291 =>	x"15000000",
		292 =>	x"16171819",
		293 =>	x"1A1B1C1D",
		294 =>	x"1E0F121F",
		295 =>	x"20191819",
		296 =>	x"210F2223",
		297 =>	x"24252627",
		298 =>	x"2819292A",
		299 =>	x"2B2C2D11",
		300 =>	x"2E2F3031",
		301 =>	x"3233342A",
		302 =>	x"35333637",
		303 =>	x"3827393A",
		304 =>	x"3B3B3B3B",
		305 =>	x"3B3B3B3B",
		306 =>	x"3B3B3B3B",
		307 =>	x"3C3D3E03",
		308 =>	x"3B3B3B3B",
		309 =>	x"3B3B3B3B",
		310 =>	x"3B3B3B3B",
		311 =>	x"3B3B3B3B",
		312 =>	x"3F404142",
		313 =>	x"4344453B",
		314 =>	x"46474849",
		315 =>	x"044A3B3B",
		316 =>	x"4B4C4D4E",
		317 =>	x"4F505152",
		318 =>	x"53545155",
		319 =>	x"56575859",
		320 =>	x"5A5B5C5D", -- IMG_16x16_car_blue
		321 =>	x"5A5B5C5D",
		322 =>	x"0000005D",
		323 =>	x"005A5E00",
		324 =>	x"5A5B5C5D",
		325 =>	x"5A5A5E5D",
		326 =>	x"005A0000",
		327 =>	x"005E5C5D",
		328 =>	x"00005E00",
		329 =>	x"0000005D",
		330 =>	x"005B5C5D",
		331 =>	x"5A5B5C5D",
		332 =>	x"00005E5D",
		333 =>	x"005A5E5F",
		334 =>	x"5C605F5D",
		335 =>	x"5A5B5C5D",
		336 =>	x"5A605B5F",
		337 =>	x"5C605F5D",
		338 =>	x"5A5B5C5D",
		339 =>	x"5A5B5E00",
		340 =>	x"5C5B5C5D",
		341 =>	x"5A5B5C5D",
		342 =>	x"5A5A0000",
		343 =>	x"005E5C5D",
		344 =>	x"00005E00",
		345 =>	x"00000000",
		346 =>	x"5A5B5C5D",
		347 =>	x"5C605B5F",
		348 =>	x"00005E5D",
		349 =>	x"005A5E5F",
		350 =>	x"5C605F5D",
		351 =>	x"5A5B5C5D",
		352 =>	x"5A5B5C5D",
		353 =>	x"5A5B5C5D",
		354 =>	x"5A5B5E5D",
		355 =>	x"005A5E00",
		356 =>	x"5A5B5E00",
		357 =>	x"00005E5D",
		358 =>	x"005A0000",
		359 =>	x"005A5C5D",
		360 =>	x"00000000",
		361 =>	x"00000000",
		362 =>	x"5A5B5C5D",
		363 =>	x"5A5B5C5D",
		364 =>	x"00000000",
		365 =>	x"005A0000",
		366 =>	x"005E5C5D",
		367 =>	x"00000000",
		368 =>	x"005A0000",
		369 =>	x"5A5A0000",
		370 =>	x"00000000",
		371 =>	x"00000000",
		372 =>	x"00000000",
		373 =>	x"00000000",
		374 =>	x"00000000",
		375 =>	x"00005E5D",
		376 =>	x"00000000",
		377 =>	x"00000000",
		378 =>	x"005A5E5D",
		379 =>	x"00000000",
		380 =>	x"00000000",
		381 =>	x"00000000",
		382 =>	x"00000000",
		383 =>	x"00000000",
		384 =>	x"5D5A5B5C", -- IMG_16x16_car_red
		385 =>	x"5D5A5B5C",
		386 =>	x"0000005D",
		387 =>	x"005A5E00",
		388 =>	x"5D5A5B5C",
		389 =>	x"5D5A5E5D",
		390 =>	x"005A0000",
		391 =>	x"00005B5C",
		392 =>	x"00005E00",
		393 =>	x"0000005D",
		394 =>	x"005A5B5C",
		395 =>	x"5D5A5B5C",
		396 =>	x"00005E5D",
		397 =>	x"005A5E5F",
		398 =>	x"5C605B5C",
		399 =>	x"5D5A5B5C",
		400 =>	x"5D605B5F",
		401 =>	x"5C605B5C",
		402 =>	x"5D5A5B5C",
		403 =>	x"5D5A5B00",
		404 =>	x"5C5A5B5C",
		405 =>	x"5D5A5B5C",
		406 =>	x"5D5A0000",
		407 =>	x"00005B5C",
		408 =>	x"00005E00",
		409 =>	x"00000000",
		410 =>	x"5D5A5B5C",
		411 =>	x"5C605B5F",
		412 =>	x"00005E5D",
		413 =>	x"005A5E5F",
		414 =>	x"5C605B5C",
		415 =>	x"5D5A5B5C",
		416 =>	x"5D5A5B5C",
		417 =>	x"5D5A5B5C",
		418 =>	x"5D5A5B5D",
		419 =>	x"005A5E00",
		420 =>	x"5D5A5B00",
		421 =>	x"00005E5D",
		422 =>	x"005A0000",
		423 =>	x"005A5E5C",
		424 =>	x"00000000",
		425 =>	x"00000000",
		426 =>	x"5D5A5B5C",
		427 =>	x"5D5A5B5C",
		428 =>	x"00000000",
		429 =>	x"005A0000",
		430 =>	x"00005B5C",
		431 =>	x"00000000",
		432 =>	x"005A0000",
		433 =>	x"5D5A0000",
		434 =>	x"00000000",
		435 =>	x"00000000",
		436 =>	x"00000000",
		437 =>	x"00000000",
		438 =>	x"00000000",
		439 =>	x"00005E5D",
		440 =>	x"00000000",
		441 =>	x"00000000",
		442 =>	x"005A5E5D",
		443 =>	x"00000000",
		444 =>	x"00000000",
		445 =>	x"00000000",
		446 =>	x"00000000",
		447 =>	x"00000000",
		448 =>	x"5C605B5F", -- IMG_16x16_flag
		449 =>	x"5C605B5F",
		450 =>	x"00000000",
		451 =>	x"00000000",
		452 =>	x"5C605B5F",
		453 =>	x"5C5A0000",
		454 =>	x"00000000",
		455 =>	x"005D5B5F",
		456 =>	x"00000000",
		457 =>	x"00000000",
		458 =>	x"5C605B5F",
		459 =>	x"5C605B5F",
		460 =>	x"0000005F",
		461 =>	x"5C605B5F",
		462 =>	x"5C605B5F",
		463 =>	x"5C5A0000",
		464 =>	x"5C605B5F",
		465 =>	x"5C5A0000",
		466 =>	x"00000000",
		467 =>	x"00000000",
		468 =>	x"00000000",
		469 =>	x"00000000",
		470 =>	x"00000000",
		471 =>	x"005D5B5F",
		472 =>	x"00000000",
		473 =>	x"00000000",
		474 =>	x"5C605B5F",
		475 =>	x"5C5A0000",
		476 =>	x"0000005F",
		477 =>	x"5C5A0000",
		478 =>	x"00000000",
		479 =>	x"00000000",
		480 =>	x"00000000",
		481 =>	x"00000000",
		482 =>	x"00000000",
		483 =>	x"00000000",
		484 =>	x"00000000",
		485 =>	x"00000000",
		486 =>	x"00000000",
		487 =>	x"005D5B5F",
		488 =>	x"00000000",
		489 =>	x"00000000",
		490 =>	x"5C605B00",
		491 =>	x"00000000",
		492 =>	x"0000005F",
		493 =>	x"5C5A0000",
		494 =>	x"00000000",
		495 =>	x"00000000",
		496 =>	x"5C5A0000",
		497 =>	x"00000000",
		498 =>	x"00000000",
		499 =>	x"00000000",
		500 =>	x"00000000",
		501 =>	x"00000000",
		502 =>	x"00000000",
		503 =>	x"5C605B5F",
		504 =>	x"00000000",
		505 =>	x"0000005F",
		506 =>	x"5C605B5F",
		507 =>	x"00000000",
		508 =>	x"00000000",
		509 =>	x"00000000",
		510 =>	x"00000000",
		511 =>	x"00000000",
		512 =>	x"00000000", -- IMG_16x16_map_element_00
		513 =>	x"00010203",
		514 =>	x"0405610A",
		515 =>	x"62636403",
		516 =>	x"00000000",
		517 =>	x"00000000",
		518 =>	x"0708090A",
		519 =>	x"0B000000",
		520 =>	x"00000000",
		521 =>	x"00000000",
		522 =>	x"00000000",
		523 =>	x"00000000",
		524 =>	x"00000000",
		525 =>	x"00000000",
		526 =>	x"00000000",
		527 =>	x"00000000",
		528 =>	x"00000000",
		529 =>	x"00000000",
		530 =>	x"00000000",
		531 =>	x"00000000",
		532 =>	x"00000000",
		533 =>	x"00000000",
		534 =>	x"00000000",
		535 =>	x"00000000",
		536 =>	x"00000000",
		537 =>	x"00000000",
		538 =>	x"00000000",
		539 =>	x"00000000",
		540 =>	x"651B662C",
		541 =>	x"67196869",
		542 =>	x"6A6B6C1B",
		543 =>	x"00000000",
		544 =>	x"1E0F121F",
		545 =>	x"20191819",
		546 =>	x"0C0D0E0F",
		547 =>	x"1011100F",
		548 =>	x"2819292A",
		549 =>	x"2B2C2D11",
		550 =>	x"16171819",
		551 =>	x"1A1B1C1D",
		552 =>	x"35333637",
		553 =>	x"3827393A",
		554 =>	x"210F2223",
		555 =>	x"24252627",
		556 =>	x"3B3B3B6D",
		557 =>	x"326E6F03",
		558 =>	x"702F3031",
		559 =>	x"3233342A",
		560 =>	x"702F713B",
		561 =>	x"3B3B3B3B",
		562 =>	x"3B3B3B3B",
		563 =>	x"3B3B3B3B",
		564 =>	x"72737475",
		565 =>	x"76777879",
		566 =>	x"777A7B7C",
		567 =>	x"3B7D7E03",
		568 =>	x"7F808182",
		569 =>	x"63838485",
		570 =>	x"86878889",
		571 =>	x"8A8B8C8D",
		572 =>	x"778E778F",
		573 =>	x"90919293",
		574 =>	x"94959697",
		575 =>	x"98999A9B",
		576 =>	x"9C9D9E5C", -- IMG_16x16_map_element_01
		577 =>	x"9C9D9E5C",
		578 =>	x"9C9D9E5C",
		579 =>	x"9C9D9F5D",
		580 =>	x"9C9D9E5C",
		581 =>	x"9C9D9E5C",
		582 =>	x"A09DA15C",
		583 =>	x"9C9D9E5C",
		584 =>	x"9C9D9EA2",
		585 =>	x"A39D9E5C",
		586 =>	x"9C9D9E5C",
		587 =>	x"9C9D9E5C",
		588 =>	x"9C9D9E5C",
		589 =>	x"9C9D9E5C",
		590 =>	x"9C9D9E5C",
		591 =>	x"9C9D9E5C",
		592 =>	x"9C9D9E5C",
		593 =>	x"9C9D9E5C",
		594 =>	x"9C9D9E5C",
		595 =>	x"9C9D9F5D",
		596 =>	x"9C9D9E5C",
		597 =>	x"9C9D9E5C",
		598 =>	x"A09DA15C",
		599 =>	x"9C9D9E5C",
		600 =>	x"9C9D9EA2",
		601 =>	x"A39D9E5C",
		602 =>	x"9C9D9E5C",
		603 =>	x"9C9D9E5C",
		604 =>	x"9C9D9E5C",
		605 =>	x"9C9D9E5C",
		606 =>	x"9C9D9E5C",
		607 =>	x"9C9D9E5C",
		608 =>	x"9C9D9E5C",
		609 =>	x"9C9D9E5C",
		610 =>	x"9C9D9E5C",
		611 =>	x"9C9D9F5D",
		612 =>	x"9C9D9E5C",
		613 =>	x"9C9D9E5C",
		614 =>	x"A09DA15C",
		615 =>	x"9C9D9E5C",
		616 =>	x"9C9D9EA2",
		617 =>	x"A39D9E5C",
		618 =>	x"9C9D9E5C",
		619 =>	x"9C9D9E5C",
		620 =>	x"9C9D9E5C",
		621 =>	x"9C9D9E5C",
		622 =>	x"9C9D9E5C",
		623 =>	x"9C9D9E5C",
		624 =>	x"9C9D9E5C",
		625 =>	x"9C9D9E5C",
		626 =>	x"9C9D9E5C",
		627 =>	x"9C9D9F5D",
		628 =>	x"9C9D9E5C",
		629 =>	x"9C9D9E5C",
		630 =>	x"A09DA15C",
		631 =>	x"9C9D9E5C",
		632 =>	x"9C9D9EA2",
		633 =>	x"A39D9E5C",
		634 =>	x"9C9D9E5C",
		635 =>	x"9C9D9E5C",
		636 =>	x"9C9D9E5C",
		637 =>	x"9C9D9E5C",
		638 =>	x"9C9D9E5C",
		639 =>	x"9C9D9E5C",
		640 =>	x"9C9D9E5C", -- IMG_16x16_map_element_02
		641 =>	x"9C9D9E5C",
		642 =>	x"9C9D9E5C",
		643 =>	x"9C9D9E5C",
		644 =>	x"9C9D9E5C",
		645 =>	x"9C9D9E5C",
		646 =>	x"9C9D9E5D",
		647 =>	x"A09D9E5C",
		648 =>	x"9C9D9E5C",
		649 =>	x"9C9DA1A2",
		650 =>	x"9C9D9E5C",
		651 =>	x"9C9D9E5C",
		652 =>	x"A39D9F5C",
		653 =>	x"9C9D9E5C",
		654 =>	x"9C9D9E5C",
		655 =>	x"9C9D9E5C",
		656 =>	x"9C9D9E5C",
		657 =>	x"9C9D9E5C",
		658 =>	x"9C9D9E5C",
		659 =>	x"9C9D9E5C",
		660 =>	x"9C9D9E5C",
		661 =>	x"9C9D9E5C",
		662 =>	x"9C9D9E5D",
		663 =>	x"A09D9E5C",
		664 =>	x"9C9D9E5C",
		665 =>	x"9C9DA1A2",
		666 =>	x"9C9D9E5C",
		667 =>	x"9C9D9E5C",
		668 =>	x"A39D9F5C",
		669 =>	x"9C9D9E5C",
		670 =>	x"9C9D9E5C",
		671 =>	x"9C9D9E5C",
		672 =>	x"9C9D9E5C",
		673 =>	x"9C9D9E5C",
		674 =>	x"9C9D9E5C",
		675 =>	x"9C9D9E5C",
		676 =>	x"9C9D9E5C",
		677 =>	x"9C9D9E5C",
		678 =>	x"9C9D9E5D",
		679 =>	x"A09D9E5C",
		680 =>	x"9C9D9E5C",
		681 =>	x"9C9DA1A2",
		682 =>	x"9C9D9E5C",
		683 =>	x"9C9D9E5C",
		684 =>	x"A39D9F5C",
		685 =>	x"9C9D9E5C",
		686 =>	x"9C9D9E5C",
		687 =>	x"9C9D9E5C",
		688 =>	x"9C9D9E5C",
		689 =>	x"9C9D9E5C",
		690 =>	x"9C9D9E5C",
		691 =>	x"9C9D9E5C",
		692 =>	x"A09D9FA2",
		693 =>	x"A09D9FA2",
		694 =>	x"A09DA45D",
		695 =>	x"A59D9E5C",
		696 =>	x"A39DA15D",
		697 =>	x"A3A6A7A8",
		698 =>	x"A99DAAA2",
		699 =>	x"A09D9FA2",
		700 =>	x"ABA6AC5D",
		701 =>	x"A39DA15D",
		702 =>	x"A39DA15D",
		703 =>	x"A39DA15D",
		704 =>	x"9C9D9E5C", -- IMG_16x16_map_element_03
		705 =>	x"9C9D9E5C",
		706 =>	x"9C9D9E5C",
		707 =>	x"9C9D9E5C",
		708 =>	x"9C9D9E5C",
		709 =>	x"9C9D9E5C",
		710 =>	x"9C9D9E5C",
		711 =>	x"9C9D9E5C",
		712 =>	x"9C9D9E5C",
		713 =>	x"9C9D9E5C",
		714 =>	x"9C9D9E5C",
		715 =>	x"9C9D9E5C",
		716 =>	x"9C9D9E5C",
		717 =>	x"9C9D9E5C",
		718 =>	x"9C9D9E5C",
		719 =>	x"9C9D9E5C",
		720 =>	x"9C9D9E5C",
		721 =>	x"9C9D9E5C",
		722 =>	x"9C9D9E5C",
		723 =>	x"9C9D9E5C",
		724 =>	x"9C9D9E5C",
		725 =>	x"9C9D9E5C",
		726 =>	x"9C9D9E5C",
		727 =>	x"9C9D9E5C",
		728 =>	x"9C9D9E5C",
		729 =>	x"9C9D9E5C",
		730 =>	x"9C9D9E5C",
		731 =>	x"9C9D9E5C",
		732 =>	x"9C9D9E5C",
		733 =>	x"9C9D9E5C",
		734 =>	x"9C9D9E5C",
		735 =>	x"9C9D9E5C",
		736 =>	x"9C9D9E5C",
		737 =>	x"9C9D9E5C",
		738 =>	x"9C9D9E5C",
		739 =>	x"9C9D9E5C",
		740 =>	x"9C9D9E5C",
		741 =>	x"9C9D9E5C",
		742 =>	x"9C9D9E5C",
		743 =>	x"9C9D9E5C",
		744 =>	x"9C9D9E5C",
		745 =>	x"9C9D9E5C",
		746 =>	x"9C9D9E5C",
		747 =>	x"9C9D9E5C",
		748 =>	x"9C9D9E5C",
		749 =>	x"9C9D9E5C",
		750 =>	x"9C9D9E5C",
		751 =>	x"9C9D9E5C",
		752 =>	x"9C9D9E5C",
		753 =>	x"9C9D9E5C",
		754 =>	x"9C9D9E5C",
		755 =>	x"9C9D9E5C",
		756 =>	x"9C9D9E5C",
		757 =>	x"9C9D9E5C",
		758 =>	x"AD9D9F5C",
		759 =>	x"9C9D9E5C",
		760 =>	x"9C9D9EA2",
		761 =>	x"A39D9FAE",
		762 =>	x"9C9D9E5C",
		763 =>	x"9C9D9E5C",
		764 =>	x"A39D9F5C",
		765 =>	x"9C9D9E5C",
		766 =>	x"9C9D9E5C",
		767 =>	x"9C9D9E5C",
		768 =>	x"9C9D9E5C", -- IMG_16x16_map_element_04
		769 =>	x"9C9D9E5C",
		770 =>	x"9C9D9E5C",
		771 =>	x"9C9D9F5D",
		772 =>	x"9C9D9E5C",
		773 =>	x"9C9D9E5C",
		774 =>	x"A09DA15C",
		775 =>	x"9C9D9E5C",
		776 =>	x"9C9D9EA2",
		777 =>	x"A39D9E5C",
		778 =>	x"9C9D9E5C",
		779 =>	x"9C9D9E5C",
		780 =>	x"9C9D9E5C",
		781 =>	x"9C9D9E5C",
		782 =>	x"9C9D9E5C",
		783 =>	x"9C9D9E5C",
		784 =>	x"9C9D9E5C",
		785 =>	x"9C9D9E5C",
		786 =>	x"9C9D9E5C",
		787 =>	x"9C9D9F5D",
		788 =>	x"9C9D9E5C",
		789 =>	x"9C9D9E5C",
		790 =>	x"A09DA15C",
		791 =>	x"9C9D9E5C",
		792 =>	x"9C9D9EA2",
		793 =>	x"A39D9E5C",
		794 =>	x"9C9D9E5C",
		795 =>	x"9C9D9E5C",
		796 =>	x"9C9D9E5C",
		797 =>	x"9C9D9E5C",
		798 =>	x"9C9D9E5C",
		799 =>	x"9C9D9E5C",
		800 =>	x"9C9D9E5C",
		801 =>	x"9C9D9E5C",
		802 =>	x"9C9D9E5C",
		803 =>	x"9C9D9F5D",
		804 =>	x"9C9D9E5C",
		805 =>	x"9C9D9E5C",
		806 =>	x"A09DA15C",
		807 =>	x"9C9D9E5C",
		808 =>	x"9C9D9EA2",
		809 =>	x"A39D9E5C",
		810 =>	x"9C9D9E5C",
		811 =>	x"9C9D9E5C",
		812 =>	x"9C9D9E5C",
		813 =>	x"9C9D9E5C",
		814 =>	x"9C9D9E5C",
		815 =>	x"9C9D9E5C",
		816 =>	x"9C9D9E5C",
		817 =>	x"9C9D9E5C",
		818 =>	x"9C9D9E5C",
		819 =>	x"9C9DAF5D",
		820 =>	x"A09D9FA2",
		821 =>	x"A09DAAB0",
		822 =>	x"B1A6A75C",
		823 =>	x"9C9D9E5C",
		824 =>	x"A3B2B3B4",
		825 =>	x"AB9D9FA2",
		826 =>	x"A09D9FA2",
		827 =>	x"A09D9FA2",
		828 =>	x"A39DA15D",
		829 =>	x"A39DA15D",
		830 =>	x"A39DA15D",
		831 =>	x"A39DA15D",
		832 =>	x"9C9D9E5C", -- IMG_16x16_map_element_05
		833 =>	x"9C9D9E5C",
		834 =>	x"9C9D9E5C",
		835 =>	x"9C9D9E5C",
		836 =>	x"9C9D9E5C",
		837 =>	x"9C9D9E5C",
		838 =>	x"9C9D9E5D",
		839 =>	x"A09D9E5C",
		840 =>	x"9C9D9E5C",
		841 =>	x"9C9DA1A2",
		842 =>	x"9C9D9E5C",
		843 =>	x"9C9D9E5C",
		844 =>	x"A39D9F5C",
		845 =>	x"9C9D9E5C",
		846 =>	x"9C9D9E5C",
		847 =>	x"9C9D9E5C",
		848 =>	x"9C9D9E5C",
		849 =>	x"9C9D9E5C",
		850 =>	x"9C9D9E5C",
		851 =>	x"9C9D9E5C",
		852 =>	x"9C9D9E5C",
		853 =>	x"9C9D9E5C",
		854 =>	x"9C9D9E5D",
		855 =>	x"A09D9E5C",
		856 =>	x"9C9D9E5C",
		857 =>	x"9C9DA1A2",
		858 =>	x"9C9D9E5C",
		859 =>	x"9C9D9E5C",
		860 =>	x"A39D9F5C",
		861 =>	x"9C9D9E5C",
		862 =>	x"9C9D9E5C",
		863 =>	x"9C9D9E5C",
		864 =>	x"9C9D9E5C",
		865 =>	x"9C9D9E5C",
		866 =>	x"9C9D9E5C",
		867 =>	x"9C9D9E5C",
		868 =>	x"9C9D9E5C",
		869 =>	x"9C9D9E5C",
		870 =>	x"9C9D9E5D",
		871 =>	x"A09D9E5C",
		872 =>	x"9C9D9E5C",
		873 =>	x"9C9DA1A2",
		874 =>	x"9C9D9E5C",
		875 =>	x"9C9D9E5C",
		876 =>	x"A39D9F5C",
		877 =>	x"9C9D9E5C",
		878 =>	x"9C9D9E5C",
		879 =>	x"9C9D9E5C",
		880 =>	x"9C9D9E5C",
		881 =>	x"9C9D9E5C",
		882 =>	x"9C9D9E5C",
		883 =>	x"9C9D9E5C",
		884 =>	x"A09D9FA2",
		885 =>	x"A09D9FA2",
		886 =>	x"A09DA45D",
		887 =>	x"A59D9E5C",
		888 =>	x"A39DA15D",
		889 =>	x"A3A6A7A8",
		890 =>	x"A99DAAA2",
		891 =>	x"A09D9FA2",
		892 =>	x"ABA6AC5D",
		893 =>	x"A39DA15D",
		894 =>	x"A39DA15D",
		895 =>	x"A39DA15D",
		896 =>	x"9C9D9E5C", -- IMG_16x16_map_element_06
		897 =>	x"9C9D9E5C",
		898 =>	x"9C9D9E5C",
		899 =>	x"9C9D9E5C",
		900 =>	x"9C9D9E5C",
		901 =>	x"9C9D9E5C",
		902 =>	x"9C9D9E5C",
		903 =>	x"9C9D9E5C",
		904 =>	x"9C9D9E5C",
		905 =>	x"9C9D9E5C",
		906 =>	x"9C9D9E5C",
		907 =>	x"9C9D9E5C",
		908 =>	x"9C9D9E5C",
		909 =>	x"9C9D9E5C",
		910 =>	x"9C9D9E5C",
		911 =>	x"9C9D9E5C",
		912 =>	x"9C9D9E5C",
		913 =>	x"9C9D9E5C",
		914 =>	x"9C9D9E5C",
		915 =>	x"9C9D9E5C",
		916 =>	x"9C9D9E5C",
		917 =>	x"9C9D9E5C",
		918 =>	x"9C9D9E5C",
		919 =>	x"9C9D9E5C",
		920 =>	x"9C9D9E5C",
		921 =>	x"9C9D9E5C",
		922 =>	x"9C9D9E5C",
		923 =>	x"9C9D9E5C",
		924 =>	x"9C9D9E5C",
		925 =>	x"9C9D9E5C",
		926 =>	x"9C9D9E5C",
		927 =>	x"9C9D9E5C",
		928 =>	x"9C9D9E5C",
		929 =>	x"9C9D9E5C",
		930 =>	x"9C9D9E5C",
		931 =>	x"9C9D9E5C",
		932 =>	x"9C9D9E5C",
		933 =>	x"9C9D9E5C",
		934 =>	x"9C9D9E5C",
		935 =>	x"9C9D9E5C",
		936 =>	x"9C9D9E5C",
		937 =>	x"9C9D9E5C",
		938 =>	x"9C9D9E5C",
		939 =>	x"9C9D9E5C",
		940 =>	x"9C9D9E5C",
		941 =>	x"9C9D9E5C",
		942 =>	x"9C9D9E5C",
		943 =>	x"9C9D9E5C",
		944 =>	x"9C9D9E5C",
		945 =>	x"9C9D9E5C",
		946 =>	x"9C9D9E5C",
		947 =>	x"9C9D9E5C",
		948 =>	x"A09D9FA2",
		949 =>	x"A09D9FA2",
		950 =>	x"A09D9F5C",
		951 =>	x"9C9D9E5C",
		952 =>	x"A39DA15D",
		953 =>	x"A39D9FA2",
		954 =>	x"A09D9FA2",
		955 =>	x"A09D9FA2",
		956 =>	x"A39DA15D",
		957 =>	x"A39DA15D",
		958 =>	x"A39DA15D",
		959 =>	x"A39DA15D",
		960 =>	x"9C9D9E5C", -- IMG_16x16_map_element_07
		961 =>	x"9C9D9E5C",
		962 =>	x"9C9D9E5C",
		963 =>	x"9C9D9F5D",
		964 =>	x"9C9D9E5C",
		965 =>	x"9C9D9E5C",
		966 =>	x"A09DA15C",
		967 =>	x"9C9D9E5C",
		968 =>	x"9C9D9EA2",
		969 =>	x"A39D9E5C",
		970 =>	x"9C9D9E5C",
		971 =>	x"9C9D9E5C",
		972 =>	x"9C9D9E5C",
		973 =>	x"9C9D9E5C",
		974 =>	x"9C9D9E5C",
		975 =>	x"9C9D9E5C",
		976 =>	x"9C9D9E5C",
		977 =>	x"9C9D9E5C",
		978 =>	x"9C9D9E5C",
		979 =>	x"9C9D9F5D",
		980 =>	x"9C9D9E5C",
		981 =>	x"9C9D9E5C",
		982 =>	x"A09DA15C",
		983 =>	x"9C9D9E5C",
		984 =>	x"9C9D9EA2",
		985 =>	x"A39D9E5C",
		986 =>	x"9C9D9E5C",
		987 =>	x"9C9D9E5C",
		988 =>	x"9C9D9E5C",
		989 =>	x"9C9D9E5C",
		990 =>	x"9C9D9E5C",
		991 =>	x"9C9D9E5C",
		992 =>	x"9C9D9E5C",
		993 =>	x"9C9D9E5C",
		994 =>	x"9C9D9E5C",
		995 =>	x"9C9D9F5D",
		996 =>	x"9C9D9E5C",
		997 =>	x"9C9D9E5C",
		998 =>	x"A09DA15C",
		999 =>	x"9C9D9E5C",
		1000 =>	x"9C9D9EA2",
		1001 =>	x"A39D9E5C",
		1002 =>	x"9C9D9E5C",
		1003 =>	x"9C9D9E5C",
		1004 =>	x"9C9D9E5C",
		1005 =>	x"9C9D9E5C",
		1006 =>	x"9C9D9E5C",
		1007 =>	x"9C9D9E5C",
		1008 =>	x"9C9D9E5C",
		1009 =>	x"9C9D9E5C",
		1010 =>	x"9C9D9E5C",
		1011 =>	x"9C9DAF5D",
		1012 =>	x"A09D9FA2",
		1013 =>	x"A09DAAB0",
		1014 =>	x"B1A6A75C",
		1015 =>	x"9C9D9E5C",
		1016 =>	x"A3B2B3B4",
		1017 =>	x"AB9D9FA2",
		1018 =>	x"A09D9FA2",
		1019 =>	x"A09D9FA2",
		1020 =>	x"A39DA15D",
		1021 =>	x"A39DA15D",
		1022 =>	x"A39DA15D",
		1023 =>	x"A39DA15D",
		1024 =>	x"9C9D9E5C", -- IMG_16x16_map_element_08
		1025 =>	x"9C9D9E5C",
		1026 =>	x"9C9D9E5C",
		1027 =>	x"9C9D9E5C",
		1028 =>	x"9C9D9E5C",
		1029 =>	x"9C9D9E5C",
		1030 =>	x"9C9D9E5D",
		1031 =>	x"A09D9E5C",
		1032 =>	x"9C9D9E5C",
		1033 =>	x"9C9DA1A2",
		1034 =>	x"9C9D9E5C",
		1035 =>	x"9C9D9E5C",
		1036 =>	x"A39D9F5C",
		1037 =>	x"9C9D9E5C",
		1038 =>	x"9C9D9E5C",
		1039 =>	x"9C9D9E5C",
		1040 =>	x"9C9D9E5C",
		1041 =>	x"9C9D9E5C",
		1042 =>	x"9C9D9E5C",
		1043 =>	x"9C9D9E5C",
		1044 =>	x"9C9D9E5C",
		1045 =>	x"9C9D9E5C",
		1046 =>	x"9C9D9E5D",
		1047 =>	x"A09D9E5C",
		1048 =>	x"9C9D9E5C",
		1049 =>	x"9C9DA1A2",
		1050 =>	x"9C9D9E5C",
		1051 =>	x"9C9D9E5C",
		1052 =>	x"A39D9F5C",
		1053 =>	x"9C9D9E5C",
		1054 =>	x"9C9D9E5C",
		1055 =>	x"9C9D9E5C",
		1056 =>	x"9C9D9E5C",
		1057 =>	x"9C9D9E5C",
		1058 =>	x"9C9D9E5C",
		1059 =>	x"9C9D9E5C",
		1060 =>	x"9C9D9E5C",
		1061 =>	x"9C9D9E5C",
		1062 =>	x"9C9D9E5D",
		1063 =>	x"A09D9E5C",
		1064 =>	x"9C9D9E5C",
		1065 =>	x"9C9DA1A2",
		1066 =>	x"9C9D9E5C",
		1067 =>	x"9C9D9E5C",
		1068 =>	x"A39D9F5C",
		1069 =>	x"9C9D9E5C",
		1070 =>	x"9C9D9E5C",
		1071 =>	x"9C9D9E5C",
		1072 =>	x"9C9D9E5C",
		1073 =>	x"9C9D9E5C",
		1074 =>	x"9C9D9E5C",
		1075 =>	x"9C9D9E5C",
		1076 =>	x"A09D9FA2",
		1077 =>	x"A09D9FA2",
		1078 =>	x"A09DA45D",
		1079 =>	x"A59D9E5C",
		1080 =>	x"A39DA15D",
		1081 =>	x"A3A6A7A8",
		1082 =>	x"A99DAAA2",
		1083 =>	x"A09D9FA2",
		1084 =>	x"ABA6AC5D",
		1085 =>	x"A39DA15D",
		1086 =>	x"A39DA15D",
		1087 =>	x"A39DA15D",
		1088 =>	x"9C9D9E5C", -- IMG_16x16_map_element_09
		1089 =>	x"9C9D9E5C",
		1090 =>	x"9C9D9E5C",
		1091 =>	x"9C9D9F5D",
		1092 =>	x"9C9D9E5C",
		1093 =>	x"9C9D9E5C",
		1094 =>	x"A09DA15D",
		1095 =>	x"A09D9E5C",
		1096 =>	x"9C9D9EA2",
		1097 =>	x"A39DA1A2",
		1098 =>	x"9C9D9E5C",
		1099 =>	x"9C9D9E5C",
		1100 =>	x"A39D9F5C",
		1101 =>	x"9C9D9E5C",
		1102 =>	x"9C9D9E5C",
		1103 =>	x"9C9D9E5C",
		1104 =>	x"9C9D9E5C",
		1105 =>	x"9C9D9E5C",
		1106 =>	x"9C9D9E5C",
		1107 =>	x"9C9D9F5D",
		1108 =>	x"9C9D9E5C",
		1109 =>	x"9C9D9E5C",
		1110 =>	x"A09DA15D",
		1111 =>	x"A09D9E5C",
		1112 =>	x"9C9D9EA2",
		1113 =>	x"A39DA1A2",
		1114 =>	x"9C9D9E5C",
		1115 =>	x"9C9D9E5C",
		1116 =>	x"A39D9F5C",
		1117 =>	x"9C9D9E5C",
		1118 =>	x"9C9D9E5C",
		1119 =>	x"9C9D9E5C",
		1120 =>	x"9C9D9E5C",
		1121 =>	x"9C9D9E5C",
		1122 =>	x"9C9D9E5C",
		1123 =>	x"9C9D9F5D",
		1124 =>	x"9C9D9E5C",
		1125 =>	x"9C9D9E5C",
		1126 =>	x"A09DA15D",
		1127 =>	x"A09D9E5C",
		1128 =>	x"9C9D9EA2",
		1129 =>	x"A39DA1A2",
		1130 =>	x"9C9D9E5C",
		1131 =>	x"9C9D9E5C",
		1132 =>	x"A39D9F5C",
		1133 =>	x"9C9D9E5C",
		1134 =>	x"9C9D9E5C",
		1135 =>	x"9C9D9E5C",
		1136 =>	x"9C9D9E5C",
		1137 =>	x"9C9D9E5C",
		1138 =>	x"9C9D9E5C",
		1139 =>	x"9C9DAF5D",
		1140 =>	x"A09D9FA2",
		1141 =>	x"A09DAAB0",
		1142 =>	x"B1A6B55D",
		1143 =>	x"A59D9E5C",
		1144 =>	x"A3B2B3B4",
		1145 =>	x"ABA6A7A8",
		1146 =>	x"A99DAAA2",
		1147 =>	x"A09D9FA2",
		1148 =>	x"ABA6AC5D",
		1149 =>	x"A39DA15D",
		1150 =>	x"A39DA15D",
		1151 =>	x"A39DA15D",
		1152 =>	x"9C9D9E5C", -- IMG_16x16_map_element_10
		1153 =>	x"9C9D9E5C",
		1154 =>	x"9C9D9E5C",
		1155 =>	x"9C9D9F5D",
		1156 =>	x"9C9D9E5C",
		1157 =>	x"9C9D9E5C",
		1158 =>	x"A09DA15C",
		1159 =>	x"9C9D9E5C",
		1160 =>	x"9C9D9EA2",
		1161 =>	x"A39D9E5C",
		1162 =>	x"9C9D9E5C",
		1163 =>	x"9C9D9E5C",
		1164 =>	x"9C9D9E5C",
		1165 =>	x"9C9D9E5C",
		1166 =>	x"9C9D9E5C",
		1167 =>	x"9C9D9E5C",
		1168 =>	x"9C9D9E5C",
		1169 =>	x"9C9D9E5C",
		1170 =>	x"9C9D9E5C",
		1171 =>	x"9C9D9F5D",
		1172 =>	x"9C9D9E5C",
		1173 =>	x"9C9D9E5C",
		1174 =>	x"A09DA15C",
		1175 =>	x"9C9D9E5C",
		1176 =>	x"9C9D9EA2",
		1177 =>	x"A39D9E5C",
		1178 =>	x"9C9D9E5C",
		1179 =>	x"9C9D9E5C",
		1180 =>	x"9C9D9E5C",
		1181 =>	x"9C9D9E5C",
		1182 =>	x"9C9D9E5C",
		1183 =>	x"9C9D9E5C",
		1184 =>	x"9C9D9E5C",
		1185 =>	x"9C9D9E5C",
		1186 =>	x"9C9D9E5C",
		1187 =>	x"9C9D9F5D",
		1188 =>	x"9C9D9E5C",
		1189 =>	x"9C9D9E5C",
		1190 =>	x"A09DA15C",
		1191 =>	x"9C9D9E5C",
		1192 =>	x"9C9D9EA2",
		1193 =>	x"A39D9E5C",
		1194 =>	x"9C9D9E5C",
		1195 =>	x"9C9D9E5C",
		1196 =>	x"9C9D9E5C",
		1197 =>	x"9C9D9E5C",
		1198 =>	x"9C9D9E5C",
		1199 =>	x"9C9D9E5C",
		1200 =>	x"9C9D9E5C",
		1201 =>	x"9C9D9E5C",
		1202 =>	x"9C9D9E5C",
		1203 =>	x"9C9DAF5D",
		1204 =>	x"A09D9FA2",
		1205 =>	x"A09DAAB0",
		1206 =>	x"B1A6A75C",
		1207 =>	x"9C9D9E5C",
		1208 =>	x"A3B2B3B4",
		1209 =>	x"AB9D9FA2",
		1210 =>	x"A09D9FA2",
		1211 =>	x"A09D9FA2",
		1212 =>	x"A39DA15D",
		1213 =>	x"A39DA15D",
		1214 =>	x"A39DA15D",
		1215 =>	x"A39DA15D",
		1216 =>	x"9C9D9E5C", -- IMG_16x16_map_element_11
		1217 =>	x"9C9D9E5C",
		1218 =>	x"9C9D9E5C",
		1219 =>	x"9C9D9E5C",
		1220 =>	x"9C9D9E5C",
		1221 =>	x"9C9D9E5C",
		1222 =>	x"9C9D9E5D",
		1223 =>	x"A09D9E5C",
		1224 =>	x"9C9D9E5C",
		1225 =>	x"9C9DA1A2",
		1226 =>	x"9C9D9E5C",
		1227 =>	x"9C9D9E5C",
		1228 =>	x"A39D9F5C",
		1229 =>	x"9C9D9E5C",
		1230 =>	x"9C9D9E5C",
		1231 =>	x"9C9D9E5C",
		1232 =>	x"9C9D9E5C",
		1233 =>	x"9C9D9E5C",
		1234 =>	x"9C9D9E5C",
		1235 =>	x"9C9D9E5C",
		1236 =>	x"9C9D9E5C",
		1237 =>	x"9C9D9E5C",
		1238 =>	x"9C9D9E5D",
		1239 =>	x"A09D9E5C",
		1240 =>	x"9C9D9E5C",
		1241 =>	x"9C9DA1A2",
		1242 =>	x"9C9D9E5C",
		1243 =>	x"9C9D9E5C",
		1244 =>	x"A39D9F5C",
		1245 =>	x"9C9D9E5C",
		1246 =>	x"9C9D9E5C",
		1247 =>	x"9C9D9E5C",
		1248 =>	x"9C9D9E5C",
		1249 =>	x"9C9D9E5C",
		1250 =>	x"9C9D9E5C",
		1251 =>	x"9C9D9E5C",
		1252 =>	x"9C9D9E5C",
		1253 =>	x"9C9D9E5C",
		1254 =>	x"9C9D9E5D",
		1255 =>	x"A09D9E5C",
		1256 =>	x"9C9D9E5C",
		1257 =>	x"9C9DA1A2",
		1258 =>	x"9C9D9E5C",
		1259 =>	x"9C9D9E5C",
		1260 =>	x"A39D9F5C",
		1261 =>	x"9C9D9E5C",
		1262 =>	x"9C9D9E5C",
		1263 =>	x"9C9D9E5C",
		1264 =>	x"9C9D9E5C",
		1265 =>	x"9C9D9E5C",
		1266 =>	x"9C9D9E5C",
		1267 =>	x"9C9D9E5C",
		1268 =>	x"9C9D9E5C",
		1269 =>	x"9C9D9E5C",
		1270 =>	x"9C9D9E5D",
		1271 =>	x"A09D9E5C",
		1272 =>	x"9C9D9E5C",
		1273 =>	x"9C9DA1A2",
		1274 =>	x"9C9D9E5C",
		1275 =>	x"9C9D9E5C",
		1276 =>	x"A39D9F5C",
		1277 =>	x"9C9D9E5C",
		1278 =>	x"9C9D9E5C",
		1279 =>	x"9C9D9E5C",
		1280 =>	x"9C9D9E5C", -- IMG_16x16_map_element_12
		1281 =>	x"9C9D9E5C",
		1282 =>	x"9C9D9E5C",
		1283 =>	x"9C9D9E5C",
		1284 =>	x"9C9D9E5C",
		1285 =>	x"9C9D9E5C",
		1286 =>	x"9C9D9E5C",
		1287 =>	x"9C9D9E5C",
		1288 =>	x"9C9D9E5C",
		1289 =>	x"9C9D9E5C",
		1290 =>	x"9C9D9E5C",
		1291 =>	x"9C9D9E5C",
		1292 =>	x"9C9D9E5C",
		1293 =>	x"9C9D9E5C",
		1294 =>	x"9C9D9E5C",
		1295 =>	x"9C9D9E5C",
		1296 =>	x"9C9D9E5C",
		1297 =>	x"9C9D9E5C",
		1298 =>	x"9C9D9E5C",
		1299 =>	x"9C9D9E5C",
		1300 =>	x"9C9D9E5C",
		1301 =>	x"9C9D9E5C",
		1302 =>	x"9C9D9E5C",
		1303 =>	x"9C9D9E5C",
		1304 =>	x"9C9D9E5C",
		1305 =>	x"9C9D9E5C",
		1306 =>	x"9C9D9E5C",
		1307 =>	x"9C9D9E5C",
		1308 =>	x"9C9D9E5C",
		1309 =>	x"9C9D9E5C",
		1310 =>	x"9C9D9E5C",
		1311 =>	x"9C9D9E5C",
		1312 =>	x"9C9D9E5C",
		1313 =>	x"9C9D9E5C",
		1314 =>	x"9C9D9E5C",
		1315 =>	x"9C9D9E5C",
		1316 =>	x"9C9D9E5C",
		1317 =>	x"9C9D9E5C",
		1318 =>	x"9C9D9E5C",
		1319 =>	x"9C9D9E5C",
		1320 =>	x"9C9D9E5C",
		1321 =>	x"9C9D9E5C",
		1322 =>	x"9C9D9E5C",
		1323 =>	x"9C9D9E5C",
		1324 =>	x"9C9D9E5C",
		1325 =>	x"9C9D9E5C",
		1326 =>	x"9C9D9E5C",
		1327 =>	x"9C9D9E5C",
		1328 =>	x"9C9D9E5C",
		1329 =>	x"9C9D9E5C",
		1330 =>	x"9C9D9E5C",
		1331 =>	x"9C9D9E5C",
		1332 =>	x"9C9D9E5C",
		1333 =>	x"9C9D9E5C",
		1334 =>	x"AD9D9F5C",
		1335 =>	x"9C9D9E5C",
		1336 =>	x"9C9D9EA2",
		1337 =>	x"A39D9FAE",
		1338 =>	x"9C9D9E5C",
		1339 =>	x"9C9D9E5C",
		1340 =>	x"A39D9F5C",
		1341 =>	x"9C9D9E5C",
		1342 =>	x"9C9D9E5C",
		1343 =>	x"9C9D9E5C",
		1344 =>	x"9C9D9E5C", -- IMG_16x16_map_element_13
		1345 =>	x"9C9D9E5C",
		1346 =>	x"9C9D9E5C",
		1347 =>	x"9C9D9E5C",
		1348 =>	x"9C9D9E5C",
		1349 =>	x"9C9D9E5C",
		1350 =>	x"9C9D9E5D",
		1351 =>	x"A09D9E5C",
		1352 =>	x"9C9D9E5C",
		1353 =>	x"9C9DA1A2",
		1354 =>	x"9C9D9E5C",
		1355 =>	x"9C9D9E5C",
		1356 =>	x"A39D9F5C",
		1357 =>	x"9C9D9E5C",
		1358 =>	x"9C9D9E5C",
		1359 =>	x"9C9D9E5C",
		1360 =>	x"9C9D9E5C",
		1361 =>	x"9C9D9E5C",
		1362 =>	x"9C9D9E5C",
		1363 =>	x"9C9D9E5C",
		1364 =>	x"9C9D9E5C",
		1365 =>	x"9C9D9E5C",
		1366 =>	x"9C9D9E5D",
		1367 =>	x"A09D9E5C",
		1368 =>	x"9C9D9E5C",
		1369 =>	x"9C9DA1A2",
		1370 =>	x"9C9D9E5C",
		1371 =>	x"9C9D9E5C",
		1372 =>	x"A39D9F5C",
		1373 =>	x"9C9D9E5C",
		1374 =>	x"9C9D9E5C",
		1375 =>	x"9C9D9E5C",
		1376 =>	x"9C9D9E5C",
		1377 =>	x"9C9D9E5C",
		1378 =>	x"9C9D9E5C",
		1379 =>	x"9C9D9E5C",
		1380 =>	x"9C9D9E5C",
		1381 =>	x"9C9D9E5C",
		1382 =>	x"9C9D9E5D",
		1383 =>	x"A09D9E5C",
		1384 =>	x"9C9D9E5C",
		1385 =>	x"9C9DA1A2",
		1386 =>	x"9C9D9E5C",
		1387 =>	x"9C9D9E5C",
		1388 =>	x"A39D9F5C",
		1389 =>	x"9C9D9E5C",
		1390 =>	x"9C9D9E5C",
		1391 =>	x"9C9D9E5C",
		1392 =>	x"9C9D9E5C",
		1393 =>	x"9C9D9E5C",
		1394 =>	x"9C9D9E5C",
		1395 =>	x"9C9D9E5C",
		1396 =>	x"9C9D9E5C",
		1397 =>	x"9C9D9E5C",
		1398 =>	x"AD9D9F5D",
		1399 =>	x"A09D9E5C",
		1400 =>	x"9C9D9EA2",
		1401 =>	x"A39DA1A2",
		1402 =>	x"9C9D9E5C",
		1403 =>	x"9C9D9E5C",
		1404 =>	x"A39D9F5C",
		1405 =>	x"9C9D9E5C",
		1406 =>	x"9C9D9E5C",
		1407 =>	x"9C9D9E5C",
		1408 =>	x"9C9D9E5C", -- IMG_16x16_map_element_14
		1409 =>	x"9C9D9E5C",
		1410 =>	x"9C9D9E5C",
		1411 =>	x"9C9D9E5C",
		1412 =>	x"9C9D9E5C",
		1413 =>	x"9C9D9E5C",
		1414 =>	x"9C9D9E5C",
		1415 =>	x"9C9D9E5C",
		1416 =>	x"9C9D9E5C",
		1417 =>	x"9C9D9E5C",
		1418 =>	x"9C9D9E5C",
		1419 =>	x"9C9D9E5C",
		1420 =>	x"9C9D9E5C",
		1421 =>	x"9C9D9E5C",
		1422 =>	x"9C9D9E5C",
		1423 =>	x"9C9D9E5C",
		1424 =>	x"9C9D9E5C",
		1425 =>	x"9C9D9E5C",
		1426 =>	x"9C9D9E5C",
		1427 =>	x"9C9D9E5C",
		1428 =>	x"9C9D9E5C",
		1429 =>	x"9C9D9E5C",
		1430 =>	x"9C9D9E5C",
		1431 =>	x"9C9D9E5C",
		1432 =>	x"9C9D9E5C",
		1433 =>	x"9C9D9E5C",
		1434 =>	x"9C9D9E5C",
		1435 =>	x"9C9D9E5C",
		1436 =>	x"9C9D9E5C",
		1437 =>	x"9C9D9E5C",
		1438 =>	x"9C9D9E5C",
		1439 =>	x"9C9D9E5C",
		1440 =>	x"9C9D9E5C",
		1441 =>	x"9C9D9E5C",
		1442 =>	x"9C9D9E5C",
		1443 =>	x"9C9D9E5C",
		1444 =>	x"9C9D9E5C",
		1445 =>	x"9C9D9E5C",
		1446 =>	x"9C9D9E5C",
		1447 =>	x"9C9D9E5C",
		1448 =>	x"9C9D9E5C",
		1449 =>	x"9C9D9E5C",
		1450 =>	x"9C9D9E5C",
		1451 =>	x"9C9D9E5C",
		1452 =>	x"9C9D9E5C",
		1453 =>	x"9C9D9E5C",
		1454 =>	x"9C9D9E5C",
		1455 =>	x"9C9D9E5C",
		1456 =>	x"9C9D9E5C",
		1457 =>	x"9C9D9E5C",
		1458 =>	x"9C9D9E5C",
		1459 =>	x"9C9D9E5C",
		1460 =>	x"A09D9FA2",
		1461 =>	x"A09D9FA2",
		1462 =>	x"A09D9F5C",
		1463 =>	x"9C9D9E5C",
		1464 =>	x"A39DA15D",
		1465 =>	x"A39D9FA2",
		1466 =>	x"A09D9FA2",
		1467 =>	x"A09D9FA2",
		1468 =>	x"A39DA15D",
		1469 =>	x"A39DA15D",
		1470 =>	x"A39DA15D",
		1471 =>	x"A39DA15D",
		1472 =>	x"9C9D9E5C", -- IMG_16x16_map_element_15
		1473 =>	x"9C9D9E5C",
		1474 =>	x"9C9D9E5C",
		1475 =>	x"9C9D9F5D",
		1476 =>	x"9C9D9E5C",
		1477 =>	x"9C9D9E5C",
		1478 =>	x"A09DA15C",
		1479 =>	x"9C9D9E5C",
		1480 =>	x"9C9D9EA2",
		1481 =>	x"A39D9E5C",
		1482 =>	x"9C9D9E5C",
		1483 =>	x"9C9D9E5C",
		1484 =>	x"9C9D9E5C",
		1485 =>	x"9C9D9E5C",
		1486 =>	x"9C9D9E5C",
		1487 =>	x"9C9D9E5C",
		1488 =>	x"9C9D9E5C",
		1489 =>	x"9C9D9E5C",
		1490 =>	x"9C9D9E5C",
		1491 =>	x"9C9D9F5D",
		1492 =>	x"9C9D9E5C",
		1493 =>	x"9C9D9E5C",
		1494 =>	x"A09DA15C",
		1495 =>	x"9C9D9E5C",
		1496 =>	x"9C9D9EA2",
		1497 =>	x"A39D9E5C",
		1498 =>	x"9C9D9E5C",
		1499 =>	x"9C9D9E5C",
		1500 =>	x"9C9D9E5C",
		1501 =>	x"9C9D9E5C",
		1502 =>	x"9C9D9E5C",
		1503 =>	x"9C9D9E5C",
		1504 =>	x"9C9D9E5C",
		1505 =>	x"9C9D9E5C",
		1506 =>	x"9C9D9E5C",
		1507 =>	x"9C9D9F5D",
		1508 =>	x"9C9D9E5C",
		1509 =>	x"9C9D9E5C",
		1510 =>	x"A09DA15C",
		1511 =>	x"9C9D9E5C",
		1512 =>	x"9C9D9EA2",
		1513 =>	x"A39D9E5C",
		1514 =>	x"9C9D9E5C",
		1515 =>	x"9C9D9E5C",
		1516 =>	x"9C9D9E5C",
		1517 =>	x"9C9D9E5C",
		1518 =>	x"9C9D9E5C",
		1519 =>	x"9C9D9E5C",
		1520 =>	x"9C9D9E5C",
		1521 =>	x"9C9D9E5C",
		1522 =>	x"9C9D9E5C",
		1523 =>	x"9C9D9F5D",
		1524 =>	x"9C9D9E5C",
		1525 =>	x"9C9D9E5C",
		1526 =>	x"A09DA15C",
		1527 =>	x"9C9D9E5C",
		1528 =>	x"9C9D9EA2",
		1529 =>	x"A39D9FAE",
		1530 =>	x"9C9D9E5C",
		1531 =>	x"9C9D9E5C",
		1532 =>	x"A39D9F5C",
		1533 =>	x"9C9D9E5C",
		1534 =>	x"9C9D9E5C",
		1535 =>	x"9C9D9E5C",
		1536 =>	x"9C9D9E5C", -- IMG_16x16_map_element_16
		1537 =>	x"9C9D9E5C",
		1538 =>	x"9C9D9E5C",
		1539 =>	x"9C9D9F5D",
		1540 =>	x"9C9D9E5C",
		1541 =>	x"9C9D9E5C",
		1542 =>	x"A09DA15D",
		1543 =>	x"A09D9E5C",
		1544 =>	x"9C9D9EA2",
		1545 =>	x"A39DA1A2",
		1546 =>	x"9C9D9E5C",
		1547 =>	x"9C9D9E5C",
		1548 =>	x"A39D9F5C",
		1549 =>	x"9C9D9E5C",
		1550 =>	x"9C9D9E5C",
		1551 =>	x"9C9D9E5C",
		1552 =>	x"9C9D9E5C",
		1553 =>	x"9C9D9E5C",
		1554 =>	x"9C9D9E5C",
		1555 =>	x"9C9D9F5D",
		1556 =>	x"9C9D9E5C",
		1557 =>	x"9C9D9E5C",
		1558 =>	x"A09DA15D",
		1559 =>	x"A09D9E5C",
		1560 =>	x"9C9D9EA2",
		1561 =>	x"A39DA1A2",
		1562 =>	x"9C9D9E5C",
		1563 =>	x"9C9D9E5C",
		1564 =>	x"A39D9F5C",
		1565 =>	x"9C9D9E5C",
		1566 =>	x"9C9D9E5C",
		1567 =>	x"9C9D9E5C",
		1568 =>	x"9C9D9E5C",
		1569 =>	x"9C9D9E5C",
		1570 =>	x"9C9D9E5C",
		1571 =>	x"9C9D9F5D",
		1572 =>	x"9C9D9E5C",
		1573 =>	x"9C9D9E5C",
		1574 =>	x"A09DA15D",
		1575 =>	x"A09D9E5C",
		1576 =>	x"9C9D9EA2",
		1577 =>	x"A39DA1A2",
		1578 =>	x"9C9D9E5C",
		1579 =>	x"9C9D9E5C",
		1580 =>	x"A39D9F5C",
		1581 =>	x"9C9D9E5C",
		1582 =>	x"9C9D9E5C",
		1583 =>	x"9C9D9E5C",
		1584 =>	x"9C9D9E5C",
		1585 =>	x"9C9D9E5C",
		1586 =>	x"9C9D9E5C",
		1587 =>	x"9C9D9F5D",
		1588 =>	x"9C9D9E5C",
		1589 =>	x"9C9D9E5C",
		1590 =>	x"A09DA15D",
		1591 =>	x"A09D9E5C",
		1592 =>	x"9C9D9EA2",
		1593 =>	x"A39DA1A2",
		1594 =>	x"9C9D9E5C",
		1595 =>	x"9C9D9E5C",
		1596 =>	x"A39D9F5C",
		1597 =>	x"9C9D9E5C",
		1598 =>	x"9C9D9E5C",
		1599 =>	x"9C9D9E5C",
		1600 =>	x"9C9D9E5C", -- IMG_16x16_map_element_17
		1601 =>	x"9C9D9E5C",
		1602 =>	x"9C9D9E5C",
		1603 =>	x"9C9D9E5C",
		1604 =>	x"9C9D9E5C",
		1605 =>	x"9C9D9E5C",
		1606 =>	x"9C9D9E5C",
		1607 =>	x"9C9D9E5C",
		1608 =>	x"9C9D9E5C",
		1609 =>	x"9C9D9E5C",
		1610 =>	x"9C9D9E5C",
		1611 =>	x"9C9D9E5C",
		1612 =>	x"9C9D9E5C",
		1613 =>	x"9C9D9E5C",
		1614 =>	x"9C9D9E5C",
		1615 =>	x"9C9D9E5C",
		1616 =>	x"9C9D9E5C",
		1617 =>	x"9C9D9E5C",
		1618 =>	x"9C9D9E5C",
		1619 =>	x"9C9D9E5C",
		1620 =>	x"9C9D9E5C",
		1621 =>	x"9C9D9E5C",
		1622 =>	x"9C9D9E5C",
		1623 =>	x"9C9D9E5C",
		1624 =>	x"9C9D9E5C",
		1625 =>	x"9C9D9E5C",
		1626 =>	x"9C9D9E5C",
		1627 =>	x"9C9D9E5C",
		1628 =>	x"9C9D9E5C",
		1629 =>	x"9C9D9E5C",
		1630 =>	x"9C9D9E5C",
		1631 =>	x"9C9D9E5C",
		1632 =>	x"9C9D9E5C",
		1633 =>	x"9C9D9E5C",
		1634 =>	x"9C9D9E5C",
		1635 =>	x"9C9D9E5C",
		1636 =>	x"9C9D9E5C",
		1637 =>	x"9C9D9E5C",
		1638 =>	x"9C9D9E5C",
		1639 =>	x"9C9D9E5C",
		1640 =>	x"9C9D9E5C",
		1641 =>	x"9C9D9E5C",
		1642 =>	x"9C9D9E5C",
		1643 =>	x"9C9D9E5C",
		1644 =>	x"9C9D9E5C",
		1645 =>	x"9C9D9E5C",
		1646 =>	x"9C9D9E5C",
		1647 =>	x"9C9D9E5C",
		1648 =>	x"9C9D9E5C",
		1649 =>	x"9C9D9E5C",
		1650 =>	x"9C9D9E5C",
		1651 =>	x"9C9D9E5C",
		1652 =>	x"A09D9FA2",
		1653 =>	x"A09D9FA2",
		1654 =>	x"A09D9F5C",
		1655 =>	x"9C9D9E5C",
		1656 =>	x"A39DA15D",
		1657 =>	x"A39D9FA2",
		1658 =>	x"A09D9FA2",
		1659 =>	x"A09D9FA2",
		1660 =>	x"A39DA15D",
		1661 =>	x"A39DA15D",
		1662 =>	x"A39DA15D",
		1663 =>	x"A39DA15D",
		1664 =>	x"9C9D9E5C", -- IMG_16x16_map_element_18
		1665 =>	x"9C9D9E5C",
		1666 =>	x"9C9D9E5C",
		1667 =>	x"9C9D9F5D",
		1668 =>	x"9C9D9E5C",
		1669 =>	x"9C9D9E5C",
		1670 =>	x"A09DA15D",
		1671 =>	x"A09D9E5C",
		1672 =>	x"9C9D9EA2",
		1673 =>	x"A39DA1A2",
		1674 =>	x"9C9D9E5C",
		1675 =>	x"9C9D9E5C",
		1676 =>	x"A39D9F5C",
		1677 =>	x"9C9D9E5C",
		1678 =>	x"9C9D9E5C",
		1679 =>	x"9C9D9E5C",
		1680 =>	x"9C9D9E5C",
		1681 =>	x"9C9D9E5C",
		1682 =>	x"9C9D9E5C",
		1683 =>	x"9C9D9F5D",
		1684 =>	x"9C9D9E5C",
		1685 =>	x"9C9D9E5C",
		1686 =>	x"A09DA15D",
		1687 =>	x"A09D9E5C",
		1688 =>	x"9C9D9EA2",
		1689 =>	x"A39DA1A2",
		1690 =>	x"9C9D9E5C",
		1691 =>	x"9C9D9E5C",
		1692 =>	x"A39D9F5C",
		1693 =>	x"9C9D9E5C",
		1694 =>	x"9C9D9E5C",
		1695 =>	x"9C9D9E5C",
		1696 =>	x"9C9D9E5C",
		1697 =>	x"9C9D9E5C",
		1698 =>	x"9C9D9E5C",
		1699 =>	x"9C9D9F5D",
		1700 =>	x"9C9D9E5C",
		1701 =>	x"9C9D9E5C",
		1702 =>	x"A09DA15D",
		1703 =>	x"A09D9E5C",
		1704 =>	x"9C9D9EA2",
		1705 =>	x"A39DA1A2",
		1706 =>	x"9C9D9E5C",
		1707 =>	x"9C9D9E5C",
		1708 =>	x"A39D9F5C",
		1709 =>	x"9C9D9E5C",
		1710 =>	x"9C9D9E5C",
		1711 =>	x"9C9D9E5C",
		1712 =>	x"9C9D9E5C",
		1713 =>	x"9C9D9E5C",
		1714 =>	x"9C9D9E5C",
		1715 =>	x"9C9DA45D",
		1716 =>	x"A09D9FA2",
		1717 =>	x"A09D9FB6",
		1718 =>	x"B7A6AC5D",
		1719 =>	x"A09D9E5C",
		1720 =>	x"A3B2B3B4",
		1721 =>	x"ABA6B8B9",
		1722 =>	x"BA9D9FA2",
		1723 =>	x"A09D9FA2",
		1724 =>	x"ABA6AC5D",
		1725 =>	x"A39DA15D",
		1726 =>	x"A39DA15D",
		1727 =>	x"A39DA15D",
		1728 =>	x"9C9D9E5C", -- IMG_16x16_map_element_19
		1729 =>	x"9C9D9E5C",
		1730 =>	x"9C9D9E5C",
		1731 =>	x"9C9D9E5C",
		1732 =>	x"9C9D9E5C",
		1733 =>	x"9C9D9E5C",
		1734 =>	x"9C9D9E5C",
		1735 =>	x"9C9D9E5C",
		1736 =>	x"9C9D9E5C",
		1737 =>	x"9C9D9E5C",
		1738 =>	x"9C9D9E5C",
		1739 =>	x"9C9D9E5C",
		1740 =>	x"9C9D9E5C",
		1741 =>	x"9C9D9E5C",
		1742 =>	x"9C9D9E5C",
		1743 =>	x"9C9D9E5C",
		1744 =>	x"9C9D9E5C",
		1745 =>	x"9C9D9E5C",
		1746 =>	x"9C9D9E5C",
		1747 =>	x"9C9D9E5C",
		1748 =>	x"9C9D9E5C",
		1749 =>	x"9C9D9E5C",
		1750 =>	x"9C9D9E5C",
		1751 =>	x"9C9D9E5C",
		1752 =>	x"9C9D9E5C",
		1753 =>	x"9C9D9E5C",
		1754 =>	x"9C9D9E5C",
		1755 =>	x"9C9D9E5C",
		1756 =>	x"9C9D9E5C",
		1757 =>	x"9C9D9E5C",
		1758 =>	x"9C9D9E5C",
		1759 =>	x"9C9D9E5C",
		1760 =>	x"9C9D9E5C",
		1761 =>	x"9C9D9E5C",
		1762 =>	x"9C9D9E5C",
		1763 =>	x"9C9D9E5C",
		1764 =>	x"9C9D9E5C",
		1765 =>	x"9C9D9E5C",
		1766 =>	x"9C9D9E5C",
		1767 =>	x"9C9D9E5C",
		1768 =>	x"9C9D9E5C",
		1769 =>	x"9C9D9E5C",
		1770 =>	x"9C9D9E5C",
		1771 =>	x"9C9D9E5C",
		1772 =>	x"9C9D9E5C",
		1773 =>	x"9C9D9E5C",
		1774 =>	x"9C9D9E5C",
		1775 =>	x"9C9D9E5C",
		1776 =>	x"9C9D9E5C",
		1777 =>	x"9C9D9E5C",
		1778 =>	x"9C9D9E5C",
		1779 =>	x"9C9D9E5C",
		1780 =>	x"9C9D9E5C",
		1781 =>	x"9C9D9E5C",
		1782 =>	x"9C9D9E5C",
		1783 =>	x"9C9D9E5C",
		1784 =>	x"9C9D9E5C",
		1785 =>	x"9C9D9E5C",
		1786 =>	x"9C9D9E5C",
		1787 =>	x"9C9D9E5C",
		1788 =>	x"9C9D9E5C",
		1789 =>	x"9C9D9E5C",
		1790 =>	x"9C9D9E5C",
		1791 =>	x"9C9D9E5C",
		1792 =>	x"9C9D9E5C", -- IMG_16x16_map_element_20
		1793 =>	x"9C9D9E5C",
		1794 =>	x"9C9D9E5C",
		1795 =>	x"9C9D9F5D",
		1796 =>	x"9C9D9E5C",
		1797 =>	x"9C9D9E5C",
		1798 =>	x"A09DA15C",
		1799 =>	x"9C9D9E5C",
		1800 =>	x"9C9D9EA2",
		1801 =>	x"A39D9E5C",
		1802 =>	x"9C9D9E5C",
		1803 =>	x"9C9D9E5C",
		1804 =>	x"9C9D9E5C",
		1805 =>	x"9C9D9E5C",
		1806 =>	x"9C9D9E5C",
		1807 =>	x"9C9D9E5C",
		1808 =>	x"9C9D9E5C",
		1809 =>	x"9C9D9E5C",
		1810 =>	x"9C9D9E5C",
		1811 =>	x"9C9D9F5D",
		1812 =>	x"9C9D9E5C",
		1813 =>	x"9C9D9E5C",
		1814 =>	x"A09DA15C",
		1815 =>	x"9C9D9E5C",
		1816 =>	x"9C9D9EA2",
		1817 =>	x"A39D9E5C",
		1818 =>	x"9C9D9E5C",
		1819 =>	x"9C9D9E5C",
		1820 =>	x"9C9D9E5C",
		1821 =>	x"9C9D9E5C",
		1822 =>	x"9C9D9E5C",
		1823 =>	x"9C9D9E5C",
		1824 =>	x"9C9D9E5C",
		1825 =>	x"9C9D9E5C",
		1826 =>	x"9C9D9E5C",
		1827 =>	x"9C9D9F5D",
		1828 =>	x"9C9D9E5C",
		1829 =>	x"9C9D9E5C",
		1830 =>	x"A09DA15C",
		1831 =>	x"9C9D9E5C",
		1832 =>	x"9C9D9EA2",
		1833 =>	x"A39D9E5C",
		1834 =>	x"9C9D9E5C",
		1835 =>	x"9C9D9E5C",
		1836 =>	x"9C9D9E5C",
		1837 =>	x"9C9D9E5C",
		1838 =>	x"9C9D9E5C",
		1839 =>	x"9C9D9E5C",
		1840 =>	x"9C9D9E5C",
		1841 =>	x"9C9D9E5C",
		1842 =>	x"9C9D9E5C",
		1843 =>	x"9C9D9F5D",
		1844 =>	x"9C9D9E5C",
		1845 =>	x"9C9D9E5C",
		1846 =>	x"A09DA15C",
		1847 =>	x"9C9D9E5C",
		1848 =>	x"9C9D9EA2",
		1849 =>	x"A39D9E5C",
		1850 =>	x"9C9D9E5C",
		1851 =>	x"9C9D9E5C",
		1852 =>	x"9C9D9E5C",
		1853 =>	x"9C9D9E5C",
		1854 =>	x"9C9D9E5C",
		1855 =>	x"9C9D9E5C",
		1856 =>	x"9C9D9E5C", -- IMG_16x16_map_element_21
		1857 =>	x"9C9D9E5C",
		1858 =>	x"9C9D9E5C",
		1859 =>	x"9C9D9E5C",
		1860 =>	x"9C9D9E5C",
		1861 =>	x"9C9D9E5C",
		1862 =>	x"9C9D9E5D",
		1863 =>	x"A09D9E5C",
		1864 =>	x"9C9D9E5C",
		1865 =>	x"9C9DA1A2",
		1866 =>	x"9C9D9E5C",
		1867 =>	x"9C9D9E5C",
		1868 =>	x"A39D9F5C",
		1869 =>	x"9C9D9E5C",
		1870 =>	x"9C9D9E5C",
		1871 =>	x"9C9D9E5C",
		1872 =>	x"9C9D9E5C",
		1873 =>	x"9C9D9E5C",
		1874 =>	x"9C9D9E5C",
		1875 =>	x"9C9D9E5C",
		1876 =>	x"9C9D9E5C",
		1877 =>	x"9C9D9E5C",
		1878 =>	x"9C9D9E5D",
		1879 =>	x"A09D9E5C",
		1880 =>	x"9C9D9E5C",
		1881 =>	x"9C9DA1A2",
		1882 =>	x"9C9D9E5C",
		1883 =>	x"9C9D9E5C",
		1884 =>	x"A39D9F5C",
		1885 =>	x"9C9D9E5C",
		1886 =>	x"9C9D9E5C",
		1887 =>	x"9C9D9E5C",
		1888 =>	x"9C9D9E5C",
		1889 =>	x"9C9D9E5C",
		1890 =>	x"9C9D9E5C",
		1891 =>	x"9C9D9E5C",
		1892 =>	x"9C9D9E5C",
		1893 =>	x"9C9D9E5C",
		1894 =>	x"9C9D9E5D",
		1895 =>	x"A09D9E5C",
		1896 =>	x"9C9D9E5C",
		1897 =>	x"9C9DA1A2",
		1898 =>	x"9C9D9E5C",
		1899 =>	x"9C9D9E5C",
		1900 =>	x"A39D9F5C",
		1901 =>	x"9C9D9E5C",
		1902 =>	x"9C9D9E5C",
		1903 =>	x"9C9D9E5C",
		1904 =>	x"9C9D9E5C",
		1905 =>	x"9C9D9E5C",
		1906 =>	x"9C9D9E5C",
		1907 =>	x"9C9D9E5C",
		1908 =>	x"9C9D9E5C",
		1909 =>	x"9C9D9E5C",
		1910 =>	x"AD9D9F5D",
		1911 =>	x"A09D9E5C",
		1912 =>	x"9C9D9EA2",
		1913 =>	x"A39DA1A2",
		1914 =>	x"9C9D9E5C",
		1915 =>	x"9C9D9E5C",
		1916 =>	x"A39D9F5C",
		1917 =>	x"9C9D9E5C",
		1918 =>	x"9C9D9E5C",
		1919 =>	x"9C9D9E5C",
		1920 =>	x"9C9D9E5C", -- IMG_16x16_map_element_22
		1921 =>	x"9C9D9E5C",
		1922 =>	x"9C9D9E5C",
		1923 =>	x"9C9D9F5D",
		1924 =>	x"9C9D9E5C",
		1925 =>	x"9C9D9E5C",
		1926 =>	x"A09DA15D",
		1927 =>	x"A09D9E5C",
		1928 =>	x"9C9D9EA2",
		1929 =>	x"A39DA1A2",
		1930 =>	x"9C9D9E5C",
		1931 =>	x"9C9D9E5C",
		1932 =>	x"A39D9F5C",
		1933 =>	x"9C9D9E5C",
		1934 =>	x"9C9D9E5C",
		1935 =>	x"9C9D9E5C",
		1936 =>	x"9C9D9E5C",
		1937 =>	x"9C9D9E5C",
		1938 =>	x"9C9D9E5C",
		1939 =>	x"9C9D9F5D",
		1940 =>	x"9C9D9E5C",
		1941 =>	x"9C9D9E5C",
		1942 =>	x"A09DA15D",
		1943 =>	x"A09D9E5C",
		1944 =>	x"9C9D9EA2",
		1945 =>	x"A39DA1A2",
		1946 =>	x"9C9D9E5C",
		1947 =>	x"9C9D9E5C",
		1948 =>	x"A39D9F5C",
		1949 =>	x"9C9D9E5C",
		1950 =>	x"9C9D9E5C",
		1951 =>	x"9C9D9E5C",
		1952 =>	x"9C9D9E5C",
		1953 =>	x"9C9D9E5C",
		1954 =>	x"9C9D9E5C",
		1955 =>	x"9C9D9F5D",
		1956 =>	x"9C9D9E5C",
		1957 =>	x"9C9D9E5C",
		1958 =>	x"A09DA15D",
		1959 =>	x"A09D9E5C",
		1960 =>	x"9C9D9EA2",
		1961 =>	x"A39DA1A2",
		1962 =>	x"9C9D9E5C",
		1963 =>	x"9C9D9E5C",
		1964 =>	x"A39D9F5C",
		1965 =>	x"9C9D9E5C",
		1966 =>	x"9C9D9E5C",
		1967 =>	x"9C9D9E5C",
		1968 =>	x"9C9D9E5C",
		1969 =>	x"9C9D9E5C",
		1970 =>	x"9C9D9E5C",
		1971 =>	x"9C9D9F5D",
		1972 =>	x"9C9D9E5C",
		1973 =>	x"9C9D9E5C",
		1974 =>	x"A09DA15D",
		1975 =>	x"A09D9E5C",
		1976 =>	x"9C9D9EA2",
		1977 =>	x"A39DA1A2",
		1978 =>	x"9C9D9E5C",
		1979 =>	x"9C9D9E5C",
		1980 =>	x"A39D9F5C",
		1981 =>	x"9C9D9E5C",
		1982 =>	x"9C9D9E5C",
		1983 =>	x"9C9D9E5C",
		1984 =>	x"9C9D9E5C", -- IMG_16x16_map_element_23
		1985 =>	x"9C9D9E5C",
		1986 =>	x"9C9D9E5C",
		1987 =>	x"9C9D9F5D",
		1988 =>	x"9C9D9E5C",
		1989 =>	x"9C9D9E5C",
		1990 =>	x"A09DA15C",
		1991 =>	x"9C9D9E5C",
		1992 =>	x"9C9D9EA2",
		1993 =>	x"A39D9E5C",
		1994 =>	x"9C9D9E5C",
		1995 =>	x"9C9D9E5C",
		1996 =>	x"9C9D9E5C",
		1997 =>	x"9C9D9E5C",
		1998 =>	x"9C9D9E5C",
		1999 =>	x"9C9D9E5C",
		2000 =>	x"9C9D9E5C",
		2001 =>	x"9C9D9E5C",
		2002 =>	x"9C9D9E5C",
		2003 =>	x"9C9D9F5D",
		2004 =>	x"9C9D9E5C",
		2005 =>	x"9C9D9E5C",
		2006 =>	x"A09DA15C",
		2007 =>	x"9C9D9E5C",
		2008 =>	x"9C9D9EA2",
		2009 =>	x"A39D9E5C",
		2010 =>	x"9C9D9E5C",
		2011 =>	x"9C9D9E5C",
		2012 =>	x"9C9D9E5C",
		2013 =>	x"9C9D9E5C",
		2014 =>	x"9C9D9E5C",
		2015 =>	x"9C9D9E5C",
		2016 =>	x"9C9D9E5C",
		2017 =>	x"9C9D9E5C",
		2018 =>	x"9C9D9E5C",
		2019 =>	x"9C9D9F5D",
		2020 =>	x"9C9D9E5C",
		2021 =>	x"9C9D9E5C",
		2022 =>	x"A09DA15C",
		2023 =>	x"9C9D9E5C",
		2024 =>	x"9C9D9EA2",
		2025 =>	x"A39D9E5C",
		2026 =>	x"9C9D9E5C",
		2027 =>	x"9C9D9E5C",
		2028 =>	x"9C9D9E5C",
		2029 =>	x"9C9D9E5C",
		2030 =>	x"9C9D9E5C",
		2031 =>	x"9C9D9E5C",
		2032 =>	x"9C9D9E5C",
		2033 =>	x"9C9D9E5C",
		2034 =>	x"9C9D9E5C",
		2035 =>	x"9C9D9F5D",
		2036 =>	x"9C9D9E5C",
		2037 =>	x"9C9D9E5C",
		2038 =>	x"A09DA15C",
		2039 =>	x"9C9D9E5C",
		2040 =>	x"9C9D9EA2",
		2041 =>	x"A39D9FAE",
		2042 =>	x"9C9D9E5C",
		2043 =>	x"9C9D9E5C",
		2044 =>	x"A39D9F5C",
		2045 =>	x"9C9D9E5C",
		2046 =>	x"9C9D9E5C",
		2047 =>	x"9C9D9E5C",
		2048 =>	x"9C9D9E5C", -- IMG_16x16_map_element_24
		2049 =>	x"9C9D9E5C",
		2050 =>	x"9C9D9E5C",
		2051 =>	x"9C9D9E5C",
		2052 =>	x"9C9D9E5C",
		2053 =>	x"9C9D9E5C",
		2054 =>	x"9C9D9E5D",
		2055 =>	x"A09D9E5C",
		2056 =>	x"9C9D9E5C",
		2057 =>	x"9C9DA1A2",
		2058 =>	x"9C9D9E5C",
		2059 =>	x"9C9D9E5C",
		2060 =>	x"A39D9F5C",
		2061 =>	x"9C9D9E5C",
		2062 =>	x"9C9D9E5C",
		2063 =>	x"9C9D9E5C",
		2064 =>	x"9C9D9E5C",
		2065 =>	x"9C9D9E5C",
		2066 =>	x"9C9D9E5C",
		2067 =>	x"9C9D9E5C",
		2068 =>	x"9C9D9E5C",
		2069 =>	x"9C9D9E5C",
		2070 =>	x"9C9D9E5D",
		2071 =>	x"A09D9E5C",
		2072 =>	x"9C9D9E5C",
		2073 =>	x"9C9DA1A2",
		2074 =>	x"9C9D9E5C",
		2075 =>	x"9C9D9E5C",
		2076 =>	x"A39D9F5C",
		2077 =>	x"9C9D9E5C",
		2078 =>	x"9C9D9E5C",
		2079 =>	x"9C9D9E5C",
		2080 =>	x"9C9D9E5C",
		2081 =>	x"9C9D9E5C",
		2082 =>	x"9C9D9E5C",
		2083 =>	x"9C9D9E5C",
		2084 =>	x"9C9D9E5C",
		2085 =>	x"9C9D9E5C",
		2086 =>	x"9C9D9E5D",
		2087 =>	x"A09D9E5C",
		2088 =>	x"9C9D9E5C",
		2089 =>	x"9C9DA1A2",
		2090 =>	x"9C9D9E5C",
		2091 =>	x"9C9D9E5C",
		2092 =>	x"A39D9F5C",
		2093 =>	x"9C9D9E5C",
		2094 =>	x"9C9D9E5C",
		2095 =>	x"9C9D9E5C",
		2096 =>	x"9C9D9E5C",
		2097 =>	x"9C9D9E5C",
		2098 =>	x"9C9D9E5C",
		2099 =>	x"9C9D9E5C",
		2100 =>	x"9C9D9E5C",
		2101 =>	x"9C9D9E5C",
		2102 =>	x"9C9D9E5D",
		2103 =>	x"A09D9E5C",
		2104 =>	x"9C9D9E5C",
		2105 =>	x"9C9DA1A2",
		2106 =>	x"9C9D9E5C",
		2107 =>	x"9C9D9E5C",
		2108 =>	x"A39D9F5C",
		2109 =>	x"9C9D9E5C",
		2110 =>	x"9C9D9E5C",
		2111 =>	x"9C9D9E5C",
		2112 =>	x"9C9D9E5C", -- IMG_16x16_map_element_25
		2113 =>	x"9C9D9E5C",
		2114 =>	x"9C9D9E5C",
		2115 =>	x"9C9D9E5C",
		2116 =>	x"9C9D9E5C",
		2117 =>	x"9C9D9E5C",
		2118 =>	x"9C9D9E5C",
		2119 =>	x"9C9D9E5C",
		2120 =>	x"9C9D9E5C",
		2121 =>	x"9C9D9E5C",
		2122 =>	x"9C9D9E5C",
		2123 =>	x"9C9D9E5C",
		2124 =>	x"9C9D9E5C",
		2125 =>	x"9C9D9E5C",
		2126 =>	x"9C9D9E5C",
		2127 =>	x"9C9D9E5C",
		2128 =>	x"9C9D9E5C",
		2129 =>	x"9C9D9E5C",
		2130 =>	x"9C9D9E5C",
		2131 =>	x"9C9D9E5C",
		2132 =>	x"9C9D9E5C",
		2133 =>	x"9C9D9E5C",
		2134 =>	x"9C9D9E5C",
		2135 =>	x"9C9D9E5C",
		2136 =>	x"9C9D9E5C",
		2137 =>	x"9C9D9E5C",
		2138 =>	x"9C9D9E5C",
		2139 =>	x"9C9D9E5C",
		2140 =>	x"9C9D9E5C",
		2141 =>	x"9C9D9E5C",
		2142 =>	x"9C9D9E5C",
		2143 =>	x"9C9D9E5C",
		2144 =>	x"9C9D9E5C",
		2145 =>	x"9C9D9E5C",
		2146 =>	x"9C9D9E5C",
		2147 =>	x"9C9D9E5C",
		2148 =>	x"9C9D9E5C",
		2149 =>	x"9C9D9E5C",
		2150 =>	x"9C9D9E5C",
		2151 =>	x"9C9D9E5C",
		2152 =>	x"9C9D9E5C",
		2153 =>	x"9C9D9E5C",
		2154 =>	x"9C9D9E5C",
		2155 =>	x"9C9D9E5C",
		2156 =>	x"9C9D9E5C",
		2157 =>	x"9C9D9E5C",
		2158 =>	x"9C9D9E5C",
		2159 =>	x"9C9D9E5C",
		2160 =>	x"9C9D9E5C",
		2161 =>	x"9C9D9E5C",
		2162 =>	x"9C9D9E5C",
		2163 =>	x"9C9D9E5C",
		2164 =>	x"9C9D9E5C",
		2165 =>	x"9C9D9E5C",
		2166 =>	x"9C9D9E5C",
		2167 =>	x"9C9D9E5C",
		2168 =>	x"9C9D9E5C",
		2169 =>	x"9C9D9E5C",
		2170 =>	x"9C9D9E5C",
		2171 =>	x"9C9D9E5C",
		2172 =>	x"9C9D9E5C",
		2173 =>	x"9C9D9E5C",
		2174 =>	x"9C9D9E5C",
		2175 =>	x"9C9D9E5C",
		2176 =>	x"00000000", -- IMG_16x16_rock
		2177 =>	x"00010203",
		2178 =>	x"0405610A",
		2179 =>	x"62636403",
		2180 =>	x"00000000",
		2181 =>	x"00000000",
		2182 =>	x"0708090A",
		2183 =>	x"0B000000",
		2184 =>	x"00000000",
		2185 =>	x"00000000",
		2186 =>	x"00000000",
		2187 =>	x"00000000",
		2188 =>	x"00000000",
		2189 =>	x"00000000",
		2190 =>	x"00000000",
		2191 =>	x"00000000",
		2192 =>	x"00000000",
		2193 =>	x"00000000",
		2194 =>	x"00000000",
		2195 =>	x"00000000",
		2196 =>	x"00000000",
		2197 =>	x"00000000",
		2198 =>	x"00000000",
		2199 =>	x"00000000",
		2200 =>	x"00000000",
		2201 =>	x"00000000",
		2202 =>	x"00000000",
		2203 =>	x"00000000",
		2204 =>	x"651B662C",
		2205 =>	x"67196869",
		2206 =>	x"BB6B6C1B",
		2207 =>	x"00000000",
		2208 =>	x"0C0D0E0F",
		2209 =>	x"1011100F",
		2210 =>	x"BC17BD0D",
		2211 =>	x"1500100F",
		2212 =>	x"16171819",
		2213 =>	x"1A1B1C1D",
		2214 =>	x"1E0F121F",
		2215 =>	x"20191819",
		2216 =>	x"210F2223",
		2217 =>	x"24252627",
		2218 =>	x"2819292A",
		2219 =>	x"2B2C2D11",
		2220 =>	x"702F3031",
		2221 =>	x"3233342A",
		2222 =>	x"35333637",
		2223 =>	x"3827393A",
		2224 =>	x"3B3B3B3B",
		2225 =>	x"3B3B3B3B",
		2226 =>	x"3B3B3B3B",
		2227 =>	x"3BBE3E03",
		2228 =>	x"3B3B3B3B",
		2229 =>	x"3B3B3B3B",
		2230 =>	x"3B3B3B3B",
		2231 =>	x"3B3B3B3B",
		2232 =>	x"BFC0C1C2",
		2233 =>	x"0044453B",
		2234 =>	x"4647C3C4",
		2235 =>	x"044A3B3B",
		2236 =>	x"C5C6C7C8",
		2237 =>	x"C9CACBCC",
		2238 =>	x"CDCECFD0",
		2239 =>	x"D1D2D3D4",
		2240 =>	x"5C605B5F", -- IMG_16x16_smoke
		2241 =>	x"5C605B5F",
		2242 =>	x"5C5A5E5F",
		2243 =>	x"5C605B5D",
		2244 =>	x"5C605B5D",
		2245 =>	x"00605B5F",
		2246 =>	x"005A0000",
		2247 =>	x"005A5E5F",
		2248 =>	x"5C605B5F",
		2249 =>	x"00605B5F",
		2250 =>	x"5C605B5F",
		2251 =>	x"005A5E5D",
		2252 =>	x"5C605B5F",
		2253 =>	x"5C5A5E5F",
		2254 =>	x"5C605B5D",
		2255 =>	x"5C605B5F",
		2256 =>	x"5C605B5F",
		2257 =>	x"5C5A5E5D",
		2258 =>	x"00605B5F",
		2259 =>	x"5C605B5D",
		2260 =>	x"5C605B5D",
		2261 =>	x"5C605B5F",
		2262 =>	x"5C5A5E00",
		2263 =>	x"5C605B5D",
		2264 =>	x"5C605B00",
		2265 =>	x"005D5B5F",
		2266 =>	x"5C5A5E5F",
		2267 =>	x"5C605B5F",
		2268 =>	x"00605B5F",
		2269 =>	x"5C605B5F",
		2270 =>	x"5C605B5F",
		2271 =>	x"5C5A5E5F",
		2272 =>	x"5C605B5F",
		2273 =>	x"5C605B5F",
		2274 =>	x"00605B5D",
		2275 =>	x"005A5E00",
		2276 =>	x"5C605B5D",
		2277 =>	x"5C605B5F",
		2278 =>	x"5C5A005F",
		2279 =>	x"5C605B5F",
		2280 =>	x"5C605B5D",
		2281 =>	x"0000005D",
		2282 =>	x"5C605B5F",
		2283 =>	x"5C605B5F",
		2284 =>	x"00005E5F",
		2285 =>	x"5C605B5F",
		2286 =>	x"5C605B5D",
		2287 =>	x"5C605B5F",
		2288 =>	x"5C5A5E5F",
		2289 =>	x"5C5A5E5F",
		2290 =>	x"5C605B5F",
		2291 =>	x"5C5A5E00",
		2292 =>	x"00605B5F",
		2293 =>	x"5C605B5D",
		2294 =>	x"005A005D",
		2295 =>	x"5C605B5F",
		2296 =>	x"005A0000",
		2297 =>	x"00005E5D",
		2298 =>	x"005A5E5D",
		2299 =>	x"00605B5F",
		2300 =>	x"00000000",
		2301 =>	x"00000000",
		2302 =>	x"005A5E00",
		2303 =>	x"00005E5D",


--			***** MAP *****


		2304 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2305 =>	x"00000140", -- z: 0 rot: 0 ptr: 320
		2306 =>	x"00000180", -- z: 0 rot: 0 ptr: 384
		2307 =>	x"00000000", -- z: 0 rot: 0 ptr: 0
		2308 =>	x"000001C0", -- z: 0 rot: 0 ptr: 448
		2309 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2310 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2311 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2312 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2313 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2314 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2315 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2316 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2317 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2318 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2319 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2320 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2321 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2322 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2323 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2324 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2325 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2326 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2327 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2328 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2329 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2330 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2331 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2332 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2333 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2334 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2335 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2336 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2337 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2338 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2339 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2340 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2341 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2342 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2343 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2344 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2345 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2346 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2347 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2348 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2349 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2350 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2351 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2352 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2353 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2354 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2355 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2356 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2357 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2358 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2359 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2360 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2361 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2362 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2363 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2364 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2365 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2366 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2367 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2368 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2369 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2370 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2371 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2372 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2373 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2374 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2375 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2377 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2378 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2379 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2380 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2381 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2382 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2383 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2384 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2385 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2386 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2387 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2388 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2389 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2390 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2391 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2392 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2393 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2394 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2395 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2396 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2397 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2398 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2399 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2400 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2401 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2402 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2403 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2404 =>	x"00000340", -- z: 0 rot: 0 ptr: 832
		2405 =>	x"00000380", -- z: 0 rot: 0 ptr: 896
		2406 =>	x"000003C0", -- z: 0 rot: 0 ptr: 960
		2407 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2408 =>	x"00000440", -- z: 0 rot: 0 ptr: 1088
		2409 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2410 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2411 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2412 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2413 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2414 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2415 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2416 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2417 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2418 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2419 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2420 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2421 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2422 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2423 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2424 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2425 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2426 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2427 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2428 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2429 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2430 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2431 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2432 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2433 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2434 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2435 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2436 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2437 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2438 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2439 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2440 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2441 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2442 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2443 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2444 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2445 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2446 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2447 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2448 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2449 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2450 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2451 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2452 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2453 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2454 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2455 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2456 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2457 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2458 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2459 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2460 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2461 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2462 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2463 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2464 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2465 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2466 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2467 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2468 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2469 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2470 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2471 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2472 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2473 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2474 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2475 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2476 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2477 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2478 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2479 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2480 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2481 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2482 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2483 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2484 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2485 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2486 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2487 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2488 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2489 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2490 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2491 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2492 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2493 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2494 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2495 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2496 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2497 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2498 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2499 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2500 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2501 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2502 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2503 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2504 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2505 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2506 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2507 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2508 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2509 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2510 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2511 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2512 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2513 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2514 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2515 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2516 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2517 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2518 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2519 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2520 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2521 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2522 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2523 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2524 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2525 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2526 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2527 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2528 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2529 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2530 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2531 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2532 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2533 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2534 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2535 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2536 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2537 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2538 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2539 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2540 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2541 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2542 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2543 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2544 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2545 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2546 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2547 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2548 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2549 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2550 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2551 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2552 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2553 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2554 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2555 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2556 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2557 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2558 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2559 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2560 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2561 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2562 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2563 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2564 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2565 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2566 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2567 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2568 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2569 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2570 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2571 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2572 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2573 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2574 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2575 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2576 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2577 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2578 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2579 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2580 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2581 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2582 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2583 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2584 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2585 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2586 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2587 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2588 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2589 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2590 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2591 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2592 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2593 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2594 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2595 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2596 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2597 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2598 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2599 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2600 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2601 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2602 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2603 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2604 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2605 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2606 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2607 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2608 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2609 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2610 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2611 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2612 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2613 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2614 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2615 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2616 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2617 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2618 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2619 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2620 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2621 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2622 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2623 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2624 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2625 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2626 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2627 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2628 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2629 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2630 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2631 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2632 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2633 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2634 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2635 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2636 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2637 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2638 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2639 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2640 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2641 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2642 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2643 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2644 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2645 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2646 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2647 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2648 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2649 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2650 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2651 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2652 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2653 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2654 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2655 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2656 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2657 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2658 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2659 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2660 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2661 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2662 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2663 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2664 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2665 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2666 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2667 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2668 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2669 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2670 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2671 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2672 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2673 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2674 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2675 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2676 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2677 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2678 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2679 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2680 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2681 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2682 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2683 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2684 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2685 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2686 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2687 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2688 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2689 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2690 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2691 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2692 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2693 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2694 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2695 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2696 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2697 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2698 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2699 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2700 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2701 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2702 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2703 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2704 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2705 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2706 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2707 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2708 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2709 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2710 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2711 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2712 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2713 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2714 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2715 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2716 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2717 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2718 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2719 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2720 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2721 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2722 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2723 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2724 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2725 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2726 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2727 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2728 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2729 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2730 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2731 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2732 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2733 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2734 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2735 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2736 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2737 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2738 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2739 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2740 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2741 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2742 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2743 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2744 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2745 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2746 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2747 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2748 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2749 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2750 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2751 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2752 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2753 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2754 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2755 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2756 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2757 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2758 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2759 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2760 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2761 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2762 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2763 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2764 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2765 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2766 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2767 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2768 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2769 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2770 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2771 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2772 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2773 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2774 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2775 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2776 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2777 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2778 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2779 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2780 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2781 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2782 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2783 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2784 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2785 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2786 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2787 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2788 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2789 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2790 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2791 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2792 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2793 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2794 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2795 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2796 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2797 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2798 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2799 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2800 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2801 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2802 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2803 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2804 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2805 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2806 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2807 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2808 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2809 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2810 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2811 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2812 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2813 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2814 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2815 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2816 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2817 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2818 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2819 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2820 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2821 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2822 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2823 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2824 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2825 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2826 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2827 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2828 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2829 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2830 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2831 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2832 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2833 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2834 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2835 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2836 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2837 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2838 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2839 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2840 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2841 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2842 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2843 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2844 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2845 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2846 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2847 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2848 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2849 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2850 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2851 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2852 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2853 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2854 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2855 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2856 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2857 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2858 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2859 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2860 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2861 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2862 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2863 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2864 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2865 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2866 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2867 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2868 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2869 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2870 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2871 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2872 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2873 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2874 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2875 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2876 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2877 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2878 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2879 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2880 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2881 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2882 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2883 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2884 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2885 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2886 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2887 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2888 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2889 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2890 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2891 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2892 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2893 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2894 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2895 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2896 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2897 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2898 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2899 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2900 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2901 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2902 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2903 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2904 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2905 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2906 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2907 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2908 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2909 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2910 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2911 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2912 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2913 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2914 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2915 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2916 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2917 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2918 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2919 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2920 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2921 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2922 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2923 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2924 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2925 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2926 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2927 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2928 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2929 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2930 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2931 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2932 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2933 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2934 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2935 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2936 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2937 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2938 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2939 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2940 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2941 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2942 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2943 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2944 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2945 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2946 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2947 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2948 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2949 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2950 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2951 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2952 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2953 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2954 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2955 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2956 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2957 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2958 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2959 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2960 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2961 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2962 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2963 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2964 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2965 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2966 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2967 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2968 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2969 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2970 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2971 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2972 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2973 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2974 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2975 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2976 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2977 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2978 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2979 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2980 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2981 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2982 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2983 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2984 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2985 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2986 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2987 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2988 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2989 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2990 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2991 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2992 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2993 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2994 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2995 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2996 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2997 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2998 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2999 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3000 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3001 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3002 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3003 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3004 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3005 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3006 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3007 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3008 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3009 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3010 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3011 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3012 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3013 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3014 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3015 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3016 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3017 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3018 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3019 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3020 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3021 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3022 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3023 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3024 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3025 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3026 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3027 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3028 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3029 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3030 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3031 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3032 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3033 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3034 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3035 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3036 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3037 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3038 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3039 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3040 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3041 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3042 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3043 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3044 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3045 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3046 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3047 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3048 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3049 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3050 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3051 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3052 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3053 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3054 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3055 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3056 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3057 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3058 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3059 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3060 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3061 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3062 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3063 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3064 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3065 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3066 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3067 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3068 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3069 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3070 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3071 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3072 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3073 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3074 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3075 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3076 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3077 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3078 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3079 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3080 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3081 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3082 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3083 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3084 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3085 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3086 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3087 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3088 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3089 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3090 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3091 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3092 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3093 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3094 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3095 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3096 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3097 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3098 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3099 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3100 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3101 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3102 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3103 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3104 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3105 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3106 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3107 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3108 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3109 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3110 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3111 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3112 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3113 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3114 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3115 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3116 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3117 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3118 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3119 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3120 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3121 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3122 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3123 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3124 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3125 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3126 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3127 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3128 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3129 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3130 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3131 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3132 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3133 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3134 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3135 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3136 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3137 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3138 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3139 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3140 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3141 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3142 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3143 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3144 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3145 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3146 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3147 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3148 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3149 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3150 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3151 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3152 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3153 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3154 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3155 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3156 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3157 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3158 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3159 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3160 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3161 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3162 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3163 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3164 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3165 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3166 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3167 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3168 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3169 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3170 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3171 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3172 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3173 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3174 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3175 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3176 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3177 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3178 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3179 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3180 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3181 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3182 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3183 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3184 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3185 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3186 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3187 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3188 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3189 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3190 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3191 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3192 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3193 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3194 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3195 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3196 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3197 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3198 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3199 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3200 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3201 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3202 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3203 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3204 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3205 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3206 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3207 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3208 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3209 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3210 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3211 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3212 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3213 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3214 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3215 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3216 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3217 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3218 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3219 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3220 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3221 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3222 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3223 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3224 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3225 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3226 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3227 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3228 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3229 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3230 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3231 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3232 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3233 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3234 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3235 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3236 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3237 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3238 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3239 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3240 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3241 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3242 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3243 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3244 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3245 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3246 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3247 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3248 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3249 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3250 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3251 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3252 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3253 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3254 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3255 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3256 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3257 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3258 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3259 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3260 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3261 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3262 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3263 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3264 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3265 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3266 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3267 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3268 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3269 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3270 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3271 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3272 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3273 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3274 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3275 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3276 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3277 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3278 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3279 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3280 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3281 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3282 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3283 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3284 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3285 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3286 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3287 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3288 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3289 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3290 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3291 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3292 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3293 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3294 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3295 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3296 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3297 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3298 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3299 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3300 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3301 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3302 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3303 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3304 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3305 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3306 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3307 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3308 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3309 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3310 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3311 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3312 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3313 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3314 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3315 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3316 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3317 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3318 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3319 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3320 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3321 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3322 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3323 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3324 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3325 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3326 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3327 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3328 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3329 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3330 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3331 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3332 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3333 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3334 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3335 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3336 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3337 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3338 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3339 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3340 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3341 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3342 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3343 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3344 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3345 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3346 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3347 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3348 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3349 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3350 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3351 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3352 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3353 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3354 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3355 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3356 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3357 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3358 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3359 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3360 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3361 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3362 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3363 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3364 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3365 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3366 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3367 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3368 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3369 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3370 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3371 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3372 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3373 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3374 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3375 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3377 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3378 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3379 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3380 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3381 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3382 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3383 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3384 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3385 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3386 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3387 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3388 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3389 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3390 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3391 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3392 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3393 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3394 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3395 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3396 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3397 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3398 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3399 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3400 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3401 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3402 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3403 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3404 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3405 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3406 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3407 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3408 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3409 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3410 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3411 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3412 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3413 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3414 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3415 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3416 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3417 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3418 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3419 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3420 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3421 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3422 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3423 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3424 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3425 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3426 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3427 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3428 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3429 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3430 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3431 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3432 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3433 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3434 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3435 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3436 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3437 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3438 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3439 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3440 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3441 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3442 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3443 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3444 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3445 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3446 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3447 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3448 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3449 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3450 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3451 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3452 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3453 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3454 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3455 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3456 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3457 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3458 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3459 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3460 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3461 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3462 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3463 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3464 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3465 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3466 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3467 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3468 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3469 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3470 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3471 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3472 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3473 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3474 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3475 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3476 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3477 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3478 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3479 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3480 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3481 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3482 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3483 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3484 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3485 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3486 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3487 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3488 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3489 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3490 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3491 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3492 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3493 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3494 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3495 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3496 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3497 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3498 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3499 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3500 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3501 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3502 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3503 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3504 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3505 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3506 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3507 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3508 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3509 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3510 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3511 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3512 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3513 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3514 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3515 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3516 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3517 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3518 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3519 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3520 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3521 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3522 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3523 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3524 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3525 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3526 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3527 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3528 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3529 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3530 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3531 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3532 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3533 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3534 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3535 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3536 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3537 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3538 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3539 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3540 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3541 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3542 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3543 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3544 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3545 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3546 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3547 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3548 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3549 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3550 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3551 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3552 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3553 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3554 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3555 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3556 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3557 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3558 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3559 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3560 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3561 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3562 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3563 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3564 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3565 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3566 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3567 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3568 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3569 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3570 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3571 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3572 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3573 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3574 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3575 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3576 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3577 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3578 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3579 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3580 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3581 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3582 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3583 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3584 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3585 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3586 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3587 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3588 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3589 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3590 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3591 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3592 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3593 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3594 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3595 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3596 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3597 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3598 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3599 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3600 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3601 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3602 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3603 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3604 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3605 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3606 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3607 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3608 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3609 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3610 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3611 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3612 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3613 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3614 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3615 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3616 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3617 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3618 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3619 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3620 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3621 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3622 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3623 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3624 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3625 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3626 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3627 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3628 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3629 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3630 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3631 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3632 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3633 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3634 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3635 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3636 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3637 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3638 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3639 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3640 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3641 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3642 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3643 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3644 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3645 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3646 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3647 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3648 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3649 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3650 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3651 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3652 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3653 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3654 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3655 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3656 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3657 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3658 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3659 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3660 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3661 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3662 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3663 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3664 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3665 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3666 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3667 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3668 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3669 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3670 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3671 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3672 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3673 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3674 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3675 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3676 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3677 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3678 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3679 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3680 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3681 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3682 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3683 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3684 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3685 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3686 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3687 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3688 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3689 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3690 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3691 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3692 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3693 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3694 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3695 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3696 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3697 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3698 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3699 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3700 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3701 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3702 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3703 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3704 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3705 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3706 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3707 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3708 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3709 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3710 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3711 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3712 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3713 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3714 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3715 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3716 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3717 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3718 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3719 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3720 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3721 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3722 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3723 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3724 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3725 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3726 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3727 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3728 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3729 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3730 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3731 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3732 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3733 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3734 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3735 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3736 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3737 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3738 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3739 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3740 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3741 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3742 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3743 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3744 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3745 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3746 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3747 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3748 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3749 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3750 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3751 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3752 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3753 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3754 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3755 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3756 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3757 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3758 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3759 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3760 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3761 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3762 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3763 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3764 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3765 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3766 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3767 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3768 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3769 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3770 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3771 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3772 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3773 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3774 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3775 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3776 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3777 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3778 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3779 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3780 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3781 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3782 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3783 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3784 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3785 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3786 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3787 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3788 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3789 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3790 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3791 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3792 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3793 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3794 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3795 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3796 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3797 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3798 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3799 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3800 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3801 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3802 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3803 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3804 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3805 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3806 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3807 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3808 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3809 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3810 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3811 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3812 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3813 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3814 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3815 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3816 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3817 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3818 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3819 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3820 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3821 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3822 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3823 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3824 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3825 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3826 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3827 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3828 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3829 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3830 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3831 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3832 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3833 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3834 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3835 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3836 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3837 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3838 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3839 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3840 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3841 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3842 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3843 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3844 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3845 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3846 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3847 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3848 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3849 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3850 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3851 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3852 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3853 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3854 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3855 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3856 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3857 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3858 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3859 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3860 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3861 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3862 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3863 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3864 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3865 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3866 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3867 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3868 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3869 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3870 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3871 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3872 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3873 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3874 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3875 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3876 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3877 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3878 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3879 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3880 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3881 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3882 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3883 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3884 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3885 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3886 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3887 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3888 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3889 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3890 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3891 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3892 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3893 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3894 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3895 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3896 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3897 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3898 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3899 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3900 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3901 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3902 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3903 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3904 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3905 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3906 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3907 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3908 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3909 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3910 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3911 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3912 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3913 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3914 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3915 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3916 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3917 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3918 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3919 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3920 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3921 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3922 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3923 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3924 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3925 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3926 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3927 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3928 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3929 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3930 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3931 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3932 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3933 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3934 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3935 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3936 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3937 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3938 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3939 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3940 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3941 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3942 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3943 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3944 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3945 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3946 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3947 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3948 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3949 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3950 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3951 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3952 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3953 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3954 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3955 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3956 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3957 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3958 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3959 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3960 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3961 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3962 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3963 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3964 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3965 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3966 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3967 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3968 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3969 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3970 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3971 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3972 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3973 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3974 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3975 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3976 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3977 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3978 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3979 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3980 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3981 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3982 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3983 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3984 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3985 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3986 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3987 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3988 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3989 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3990 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3991 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3992 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3993 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3994 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3995 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3996 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3997 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3998 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		3999 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4000 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4001 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4002 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4003 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4004 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4005 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4006 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4007 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4008 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4009 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4010 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4011 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4012 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4013 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4014 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4015 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4016 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4017 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4018 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4019 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4020 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4021 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4022 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4023 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4024 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4025 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4026 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4027 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4028 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4029 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4030 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4031 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4032 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4033 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4034 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4035 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4036 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4037 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4038 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4039 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4040 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4041 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4042 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4043 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4044 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4045 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4046 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4047 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4048 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4049 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4050 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4051 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4052 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4053 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4054 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4055 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4056 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4057 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4058 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4059 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4060 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4061 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4062 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4063 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4064 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4065 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4066 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4067 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4068 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4069 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4070 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4071 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4072 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4073 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4074 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4075 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4076 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4077 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4078 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4079 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4080 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4081 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4082 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4083 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4084 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4085 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4086 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4087 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4088 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4089 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4090 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4091 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4092 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4093 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4094 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4095 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4096 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4097 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4098 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4099 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4100 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4101 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4102 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4103 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4104 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4105 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4106 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4107 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4108 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4109 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4110 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4111 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4112 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4113 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4114 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4115 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4116 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4117 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4118 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4119 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4120 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4121 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4122 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4123 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4124 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4125 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4126 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4127 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4128 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4129 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4130 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4131 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4132 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4133 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4134 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4135 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4136 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4137 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4138 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4139 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4140 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4141 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4142 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4143 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4144 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4145 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4146 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4147 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4148 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4149 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4150 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4151 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4152 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4153 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4154 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4155 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4156 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4157 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4158 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4159 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4160 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4161 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4162 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4163 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4164 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4165 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4166 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4167 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4168 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4169 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4170 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4171 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4172 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4173 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4174 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4175 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4176 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4177 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4178 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4179 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4180 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4181 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4182 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4183 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4184 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4185 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4186 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4187 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4188 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4189 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4190 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4191 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4192 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4193 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4194 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4195 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4196 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4197 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4198 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4199 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4200 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4201 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4202 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4203 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4204 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4205 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4206 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4207 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4208 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4209 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4210 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4211 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4212 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4213 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4214 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4215 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4216 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4217 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4218 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4219 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4220 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4221 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4222 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4223 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4224 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4225 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4226 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4227 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4228 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4229 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4230 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4231 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4232 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4233 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4234 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4235 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4236 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4237 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4238 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4239 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4240 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4241 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4242 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4243 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4244 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4245 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4246 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4247 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4248 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4249 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4250 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4251 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4252 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4253 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4254 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4255 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4256 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4257 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4258 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4259 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4260 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4261 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4262 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4263 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4264 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4265 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4266 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4267 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4268 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4269 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4270 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4271 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4272 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4273 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4274 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4275 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4276 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4277 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4278 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4279 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4280 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4281 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4282 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4283 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4284 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4285 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4286 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4287 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4288 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4289 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4290 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4291 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4292 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4293 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4294 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4295 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4296 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4297 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4298 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4299 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4300 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4301 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4302 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4303 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4304 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4305 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4306 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4307 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4308 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4309 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4310 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4311 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4312 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4313 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4314 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4315 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4316 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4317 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4318 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4319 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4320 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4321 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4322 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4323 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4324 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4325 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4326 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4327 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4328 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4329 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4330 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4331 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4332 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4333 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4334 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4335 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4336 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4337 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4338 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4339 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4340 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4341 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4342 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4343 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4344 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4345 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4346 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4347 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4348 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4349 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4350 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4351 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4352 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4353 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4354 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4355 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4356 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4357 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4358 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4359 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4360 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4361 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4362 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4363 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4364 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4365 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4366 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4367 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4368 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4369 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4370 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4371 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4372 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4373 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4374 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4375 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4377 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4378 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4379 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4380 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4381 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4382 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4383 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4384 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4385 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4386 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4387 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4388 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4389 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4390 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4391 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4392 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4393 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4394 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4395 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4396 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4397 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4398 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4399 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4400 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4401 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4402 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4403 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4404 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4405 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4406 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4407 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4408 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4409 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4410 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4411 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4412 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4413 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4414 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4415 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4416 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4417 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4418 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4419 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4420 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4421 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4422 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4423 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4424 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4425 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4426 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4427 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4428 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4429 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4430 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4431 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4432 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4433 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4434 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4435 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4436 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4437 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4438 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4439 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4440 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4441 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4442 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4443 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4444 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4445 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4446 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4447 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4448 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4449 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4450 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4451 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4452 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4453 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4454 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4455 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4456 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4457 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4458 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4459 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4460 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4461 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4462 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4463 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4464 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4465 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4466 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4467 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4468 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4469 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4470 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4471 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4472 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4473 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4474 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4475 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4476 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4477 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4478 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4479 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4480 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4481 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4482 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4483 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4484 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4485 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4486 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4487 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4488 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4489 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4490 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4491 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4492 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4493 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4494 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4495 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4496 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4497 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4498 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4499 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4500 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4501 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4502 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4503 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4504 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4505 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4506 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4507 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4508 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4509 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4510 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4511 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4512 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4513 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4514 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4515 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4516 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4517 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4518 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4519 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4520 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4521 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4522 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4523 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4524 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4525 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4526 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4527 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4528 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4529 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4530 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4531 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4532 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4533 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4534 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4535 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4536 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4537 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4538 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4539 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4540 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4541 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4542 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4543 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4544 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4545 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4546 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4547 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4548 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4549 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4550 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4551 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4552 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4553 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4554 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4555 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4556 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4557 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4558 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4559 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4560 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4561 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4562 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4563 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4564 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4565 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4566 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4567 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4568 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4569 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4570 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4571 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4572 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4573 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4574 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4575 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4576 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4577 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4578 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4579 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4580 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4581 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4582 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4583 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4584 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4585 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4586 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4587 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4588 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4589 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4590 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4591 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4592 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4593 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4594 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4595 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4596 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4597 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4598 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4599 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4600 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4601 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4602 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4603 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4604 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4605 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4606 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4607 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4608 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4609 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4610 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4611 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4612 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4613 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4614 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4615 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4616 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4617 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4618 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4619 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4620 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4621 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4622 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4623 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4624 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4625 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4626 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4627 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4628 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4629 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4630 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4631 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4632 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4633 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4634 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4635 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4636 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4637 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4638 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4639 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4640 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4641 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4642 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4643 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4644 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4645 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4646 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4647 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4648 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4649 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4650 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4651 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4652 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4653 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4654 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4655 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4656 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4657 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4658 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4659 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4660 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4661 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4662 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4663 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4664 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4665 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4666 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4667 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4668 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4669 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4670 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4671 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4672 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4673 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4674 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4675 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4676 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4677 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4678 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4679 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4680 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4681 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4682 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4683 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4684 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4685 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4686 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4687 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4688 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4689 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4690 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4691 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4692 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4693 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4694 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4695 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4696 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4697 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4698 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4699 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4700 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4701 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4702 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4703 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4704 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4705 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4706 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4707 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4708 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4709 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4710 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4711 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4712 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4713 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4714 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4715 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4716 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4717 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4718 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4719 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4720 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4721 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4722 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4723 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4724 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4725 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4726 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4727 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4728 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4729 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4730 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4731 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4732 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4733 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4734 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4735 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4736 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4737 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4738 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4739 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4740 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4741 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4742 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4743 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4744 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4745 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4746 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4747 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4748 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4749 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4750 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4751 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4752 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4753 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4754 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4755 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4756 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4757 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4758 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4759 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4760 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4761 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4762 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4763 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4764 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4765 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4766 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4767 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4768 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4769 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4770 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4771 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4772 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4773 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4774 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4775 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4776 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4777 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4778 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4779 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4780 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4781 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4782 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4783 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4784 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4785 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4786 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4787 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4788 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4789 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4790 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4791 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4792 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4793 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4794 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4795 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4796 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4797 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4798 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4799 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4800 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4801 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4802 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4803 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4804 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4805 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4806 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4807 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4808 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4809 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4810 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4811 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4812 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4813 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4814 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4815 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4816 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4817 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4818 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4819 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4820 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4821 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4822 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4823 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4824 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4825 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4826 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4827 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4828 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4829 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4830 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4831 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4832 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4833 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4834 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4835 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4836 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4837 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4838 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4839 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4840 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4841 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4842 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4843 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4844 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4845 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4846 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4847 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4848 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4849 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4850 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4851 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4852 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4853 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4854 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4855 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4856 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4857 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4858 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4859 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4860 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4861 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4862 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4863 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4864 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4865 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4866 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4867 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4868 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4869 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4870 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4871 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4872 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4873 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4874 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4875 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4876 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4877 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4878 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4879 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4880 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4881 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4882 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4883 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4884 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4885 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4886 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4887 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4888 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4889 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4890 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4891 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4892 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4893 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4894 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4895 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4896 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4897 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4898 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4899 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4900 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4901 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4902 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4903 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4904 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4905 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4906 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4907 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4908 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4909 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4910 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4911 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4912 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4913 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4914 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4915 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4916 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4917 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4918 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4919 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4920 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4921 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4922 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4923 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4924 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4925 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4926 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4927 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4928 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4929 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4930 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4931 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4932 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4933 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4934 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4935 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4936 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4937 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4938 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4939 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4940 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4941 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4942 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4943 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4944 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4945 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4946 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4947 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4948 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4949 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4950 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4951 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4952 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4953 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4954 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4955 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4956 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4957 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4958 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4959 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4960 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4961 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4962 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4963 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4964 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4965 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4966 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4967 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4968 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4969 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4970 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4971 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4972 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4973 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4974 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4975 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4976 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4977 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4978 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4979 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4980 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4981 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4982 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4983 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4984 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4985 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4986 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4987 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4988 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4989 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4990 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4991 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4992 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4993 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4994 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4995 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4996 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4997 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4998 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		4999 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5000 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5001 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5002 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5003 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5004 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5005 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5006 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5007 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5008 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5009 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5010 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5011 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5012 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5013 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5014 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5015 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5016 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5017 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5018 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5019 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5020 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5021 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5022 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5023 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5024 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5025 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5026 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5027 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5028 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5029 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5030 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5031 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5032 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5033 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5034 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5035 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5036 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5037 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5038 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5039 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5040 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5041 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5042 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5043 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5044 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5045 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5046 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5047 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5048 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5049 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5050 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5051 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5052 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5053 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5054 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5055 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5056 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5057 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5058 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5059 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5060 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5061 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5062 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5063 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5064 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5065 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5066 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5067 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5068 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5069 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5070 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5071 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5072 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5073 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5074 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5075 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5076 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5077 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5078 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5079 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5080 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5081 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5082 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5083 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5084 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5085 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5086 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5087 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5088 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5089 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5090 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5091 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5092 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5093 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5094 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5095 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5096 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5097 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5098 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5099 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5100 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5101 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5102 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5103 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5104 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5105 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5106 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5107 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5108 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5109 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5110 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5111 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5112 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5113 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5114 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5115 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5116 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5117 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5118 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5119 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5120 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5121 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5122 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5123 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5124 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5125 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5126 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5127 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5128 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5129 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5130 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5131 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5132 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5133 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5134 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5135 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5136 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5137 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5138 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5139 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5140 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5141 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5142 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5143 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5144 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5145 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5146 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5147 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5148 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5149 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5150 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5151 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5152 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5153 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5154 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5155 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5156 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5157 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5158 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5159 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5160 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5161 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5162 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5163 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5164 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5165 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5166 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5167 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5168 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5169 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5170 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5171 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5172 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5173 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5174 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5175 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5176 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5177 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5178 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5179 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5180 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5181 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5182 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5183 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5184 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5185 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5186 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5187 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5188 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5189 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5190 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5191 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5192 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5193 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5194 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5195 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5196 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5197 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5198 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5199 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5200 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5201 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5202 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5203 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5204 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5205 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5206 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5207 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5208 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5209 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5210 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5211 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5212 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5213 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5214 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5215 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5216 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5217 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5218 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5219 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5220 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5221 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5222 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5223 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5224 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5225 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5226 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5227 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5228 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5229 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5230 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5231 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5232 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5233 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5234 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5235 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5236 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5237 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5238 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5239 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5240 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5241 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5242 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5243 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5244 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5245 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5246 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5247 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5248 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5249 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5250 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5251 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5252 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5253 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5254 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5255 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5256 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5257 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5258 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5259 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5260 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5261 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5262 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5263 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5264 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5265 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5266 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5267 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5268 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5269 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5270 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5271 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5272 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5273 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5274 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5275 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5276 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5277 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5278 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5279 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5280 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5281 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5282 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5283 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5284 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5285 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5286 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5287 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5288 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5289 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5290 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5291 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5292 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5293 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5294 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5295 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5296 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5297 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5298 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5299 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5300 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5301 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5302 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5303 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5304 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5305 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5306 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5307 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5308 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5309 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5310 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5311 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5312 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5313 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5314 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5315 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5316 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5317 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5318 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5319 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5320 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5321 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5322 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5323 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5324 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5325 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5326 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5327 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5328 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5329 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5330 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5331 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5332 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5333 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5334 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5335 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5336 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5337 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5338 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5339 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5340 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5341 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5342 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5343 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5344 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5345 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5346 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5347 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5348 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5349 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5350 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5351 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5352 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5353 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5354 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5355 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5356 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5357 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5358 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5359 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5360 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5361 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5362 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5363 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5364 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5365 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5366 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5367 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5368 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5369 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5370 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5371 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5372 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5373 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5374 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5375 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5377 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5378 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5379 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5380 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5381 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5382 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5383 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5384 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5385 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5386 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5387 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5388 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5389 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5390 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5391 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5392 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5393 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5394 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5395 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5396 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5397 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5398 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5399 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5400 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5401 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5402 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5403 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5404 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5405 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5406 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5407 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5408 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5409 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5410 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5411 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5412 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5413 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5414 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5415 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5416 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5417 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5418 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5419 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5420 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5421 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5422 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5423 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5424 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5425 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5426 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5427 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5428 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5429 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5430 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5431 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5432 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5433 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5434 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5435 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5436 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5437 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5438 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5439 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5440 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5441 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5442 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5443 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5444 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5445 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5446 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5447 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5448 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5449 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5450 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5451 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5452 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5453 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5454 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5455 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5456 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5457 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5458 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5459 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5460 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5461 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5462 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5463 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5464 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5465 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5466 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5467 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5468 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5469 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5470 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5471 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5472 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5473 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5474 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5475 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5476 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5477 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5478 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5479 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5480 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5481 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5482 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5483 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5484 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5485 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5486 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5487 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5488 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5489 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5490 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5491 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5492 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5493 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5494 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5495 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5496 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5497 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5498 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5499 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5500 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5501 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5502 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5503 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5504 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5505 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5506 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5507 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5508 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5509 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5510 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5511 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5512 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5513 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5514 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5515 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5516 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5517 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5518 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5519 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5520 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5521 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5522 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5523 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5524 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5525 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5526 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5527 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5528 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5529 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5530 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5531 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5532 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5533 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5534 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5535 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5536 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5537 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5538 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5539 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5540 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5541 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5542 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5543 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5544 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5545 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5546 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5547 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5548 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5549 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5550 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5551 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5552 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5553 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5554 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5555 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5556 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5557 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5558 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5559 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5560 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5561 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5562 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5563 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5564 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5565 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5566 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5567 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5568 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5569 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5570 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5571 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5572 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5573 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5574 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5575 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5576 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5577 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5578 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5579 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5580 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5581 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5582 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5583 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5584 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5585 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5586 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5587 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5588 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5589 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5590 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5591 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5592 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5593 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5594 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5595 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5596 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5597 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5598 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5599 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5600 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5601 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5602 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5603 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5604 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5605 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5606 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5607 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5608 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5609 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5610 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5611 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5612 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5613 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5614 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5615 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5616 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5617 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5618 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5619 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5620 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5621 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5622 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5623 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5624 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5625 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5626 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5627 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5628 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5629 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5630 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5631 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5632 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5633 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5634 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5635 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5636 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5637 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5638 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5639 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5640 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5641 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5642 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5643 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5644 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5645 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5646 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5647 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5648 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5649 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5650 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5651 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5652 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5653 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5654 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5655 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5656 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5657 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5658 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5659 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5660 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5661 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5662 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5663 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5664 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5665 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5666 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5667 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5668 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5669 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5670 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5671 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5672 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5673 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5674 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5675 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5676 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5677 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5678 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5679 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5680 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5681 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5682 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5683 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5684 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5685 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5686 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5687 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5688 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5689 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5690 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5691 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5692 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5693 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5694 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5695 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5696 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5697 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5698 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5699 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5700 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5701 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5702 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5703 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5704 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5705 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5706 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5707 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5708 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5709 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5710 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5711 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5712 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5713 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5714 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5715 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5716 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5717 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5718 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5719 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5720 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5721 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5722 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5723 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5724 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5725 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5726 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5727 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5728 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5729 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5730 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5731 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5732 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5733 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5734 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5735 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5736 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5737 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5738 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5739 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5740 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5741 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5742 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5743 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5744 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5745 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5746 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5747 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5748 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5749 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5750 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5751 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5752 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5753 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5754 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5755 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5756 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5757 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5758 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5759 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5760 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5761 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5762 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5763 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5764 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5765 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5766 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5767 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5768 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5769 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5770 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5771 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5772 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5773 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5774 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5775 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5776 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5777 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5778 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5779 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5780 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5781 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5782 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5783 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5784 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5785 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5786 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5787 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5788 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5789 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5790 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5791 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5792 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5793 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5794 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5795 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5796 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5797 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5798 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5799 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5800 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5801 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5802 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5803 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5804 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5805 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5806 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5807 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5808 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5809 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5810 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5811 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5812 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5813 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5814 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5815 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5816 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5817 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5818 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5819 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5820 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5821 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5822 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5823 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5824 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5825 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5826 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5827 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5828 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5829 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5830 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5831 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5832 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5833 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5834 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5835 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5836 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5837 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5838 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5839 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5840 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5841 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5842 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5843 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5844 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5845 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5846 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5847 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5848 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5849 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5850 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5851 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5852 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5853 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5854 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5855 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5856 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5857 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5858 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5859 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5860 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5861 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5862 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5863 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5864 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5865 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5866 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5867 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5868 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5869 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5870 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5871 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5872 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5873 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5874 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5875 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5876 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5877 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5878 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5879 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5880 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5881 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5882 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5883 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5884 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5885 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5886 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5887 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5888 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5889 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5890 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5891 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5892 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5893 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5894 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5895 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5896 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5897 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5898 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5899 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5900 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5901 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5902 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5903 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5904 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5905 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5906 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5907 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5908 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5909 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5910 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5911 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5912 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5913 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5914 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5915 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5916 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5917 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5918 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5919 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5920 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5921 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5922 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5923 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5924 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5925 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5926 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5927 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5928 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5929 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5930 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5931 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5932 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5933 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5934 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5935 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5936 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5937 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5938 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5939 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5940 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5941 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5942 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5943 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5944 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5945 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5946 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5947 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5948 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5949 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5950 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5951 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5952 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5953 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5954 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5955 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5956 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5957 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5958 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5959 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5960 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5961 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5962 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5963 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5964 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5965 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5966 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5967 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5968 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5969 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5970 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5971 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5972 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5973 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5974 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5975 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5976 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5977 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5978 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5979 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5980 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5981 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5982 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5983 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5984 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5985 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5986 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5987 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5988 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5989 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5990 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5991 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5992 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5993 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5994 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5995 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5996 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5997 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5998 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		5999 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6000 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6001 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6002 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6003 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6004 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6005 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6006 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6007 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6008 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6009 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6010 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6011 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6012 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6013 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6014 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6015 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6016 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6017 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6018 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6019 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6020 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6021 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6022 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6023 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6024 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6025 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6026 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6027 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6028 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6029 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6030 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6031 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6032 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6033 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6034 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6035 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6036 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6037 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6038 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6039 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6040 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6041 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6042 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6043 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6044 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6045 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6046 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6047 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6048 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6049 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6050 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6051 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6052 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6053 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6054 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6055 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6056 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6057 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6058 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6059 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6060 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6061 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6062 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6063 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6064 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6065 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6066 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6067 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6068 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6069 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6070 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6071 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6072 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6073 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6074 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6075 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6076 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6077 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6078 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6079 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6080 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6081 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6082 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6083 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6084 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6085 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6086 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6087 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6088 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6089 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6090 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6091 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6092 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6093 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6094 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6095 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6096 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6097 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6098 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6099 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6100 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6101 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6102 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6103 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6104 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6105 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6106 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6107 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6108 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6109 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6110 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6111 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6112 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6113 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6114 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6115 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6116 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6117 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6118 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6119 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6120 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6121 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6122 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6123 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6124 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6125 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6126 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6127 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6128 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6129 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6130 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6131 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6132 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6133 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6134 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6135 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6136 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6137 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6138 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6139 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6140 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6141 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6142 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6143 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6144 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6145 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6146 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6147 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6148 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6149 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6150 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6151 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6152 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6153 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6154 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6155 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6156 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6157 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6158 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6159 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6160 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6161 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6162 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6163 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6164 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6165 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6166 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6167 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6168 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6169 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6170 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6171 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6172 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6173 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6174 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6175 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6176 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6177 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6178 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6179 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6180 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6181 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6182 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6183 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6184 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6185 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6186 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6187 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6188 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6189 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6190 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6191 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6192 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6193 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6194 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6195 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6196 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6197 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6198 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6199 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6200 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6201 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6202 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6203 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6204 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6205 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6206 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6207 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6208 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6209 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6210 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6211 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6212 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6213 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6214 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6215 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6216 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6217 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6218 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6219 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6220 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6221 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6222 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6223 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6224 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6225 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6226 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6227 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6228 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6229 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6230 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6231 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6232 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6233 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6234 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6235 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6236 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6237 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6238 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6239 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6240 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6241 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6242 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6243 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6244 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6245 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6246 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6247 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6248 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6249 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6250 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6251 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6252 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6253 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6254 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6255 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6256 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6257 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6258 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6259 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6260 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6261 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6262 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6263 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6264 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6265 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6266 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6267 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6268 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6269 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6270 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6271 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6272 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6273 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6274 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6275 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6276 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6277 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6278 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6279 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6280 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6281 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6282 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6283 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6284 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6285 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6286 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6287 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6288 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6289 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6290 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6291 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6292 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6293 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6294 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6295 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6296 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6297 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6298 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6299 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6300 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6301 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6302 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6303 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6304 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6305 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6306 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6307 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6308 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6309 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6310 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6311 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6312 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6313 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6314 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6315 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6316 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6317 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6318 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6319 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6320 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6321 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6322 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6323 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6324 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6325 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6326 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6327 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6328 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6329 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6330 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6331 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6332 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6333 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6334 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6335 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6336 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6337 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6338 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6339 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6340 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6341 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6342 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6343 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6344 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6345 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6346 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6347 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6348 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6349 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6350 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6351 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6352 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6353 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6354 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6355 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6356 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6357 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6358 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6359 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6360 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6361 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6362 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6363 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6364 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6365 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6366 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6367 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6368 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6369 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6370 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6371 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6372 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6373 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6374 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6375 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6377 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6378 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6379 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6380 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6381 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6382 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6383 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6384 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6385 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6386 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6387 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6388 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6389 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6390 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6391 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6392 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6393 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6394 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6395 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6396 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6397 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6398 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6399 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6400 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6401 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6402 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6403 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6404 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6405 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6406 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6407 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6408 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6409 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6410 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6411 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6412 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6413 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6414 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6415 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6416 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6417 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6418 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6419 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6420 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6421 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6422 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6423 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6424 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6425 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6426 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6427 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6428 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6429 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6430 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6431 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6432 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6433 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6434 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6435 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6436 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6437 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6438 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6439 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6440 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6441 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6442 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6443 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6444 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6445 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6446 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6447 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6448 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6449 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6450 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6451 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6452 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6453 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6454 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6455 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6456 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6457 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6458 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6459 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6460 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6461 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6462 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6463 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6464 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6465 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6466 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6467 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6468 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6469 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6470 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6471 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6472 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6473 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6474 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6475 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6476 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6477 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6478 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6479 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6480 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6481 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6482 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6483 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6484 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6485 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6486 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6487 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6488 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6489 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6490 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6491 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6492 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6493 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6494 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6495 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6496 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6497 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6498 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6499 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6500 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6501 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6502 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6503 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6504 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6505 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6506 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6507 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6508 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6509 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6510 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6511 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6512 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6513 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6514 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6515 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6516 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6517 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6518 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6519 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6520 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6521 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6522 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6523 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6524 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6525 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6526 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6527 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6528 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6529 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6530 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6531 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6532 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6533 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6534 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6535 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6536 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6537 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6538 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6539 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6540 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6541 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6542 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6543 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6544 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6545 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6546 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6547 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6548 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6549 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6550 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6551 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6552 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6553 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6554 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6555 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6556 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6557 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6558 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6559 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6560 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6561 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6562 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6563 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6564 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6565 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6566 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6567 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6568 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6569 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6570 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6571 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6572 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6573 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6574 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6575 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6576 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6577 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6578 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6579 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6580 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6581 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6582 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6583 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6584 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6585 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6586 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6587 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6588 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6589 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6590 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6591 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6592 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6593 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6594 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6595 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6596 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6597 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6598 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6599 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6600 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6601 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6602 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6603 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6604 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6605 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6606 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6607 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6608 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6609 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6610 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6611 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6612 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6613 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6614 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6615 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6616 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6617 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6618 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6619 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6620 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6621 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6622 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6623 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6624 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6625 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6626 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6627 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6628 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6629 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6630 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6631 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6632 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6633 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6634 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6635 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6636 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6637 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6638 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6639 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6640 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6641 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6642 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6643 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6644 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6645 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6646 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6647 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6648 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6649 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6650 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6651 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6652 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6653 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6654 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6655 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6656 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6657 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6658 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6659 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6660 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6661 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6662 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6663 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6664 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6665 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6666 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6667 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6668 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6669 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6670 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6671 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6672 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6673 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6674 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6675 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6676 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6677 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6678 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6679 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6680 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6681 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6682 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6683 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6684 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6685 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6686 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6687 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6688 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6689 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6690 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6691 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6692 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6693 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6694 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6695 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6696 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6697 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6698 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6699 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6700 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6701 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6702 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6703 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6704 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6705 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6706 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6707 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6708 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6709 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6710 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6711 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6712 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6713 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6714 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6715 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6716 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6717 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6718 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6719 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6720 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6721 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6722 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6723 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6724 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6725 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6726 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6727 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6728 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6729 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6730 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6731 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6732 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6733 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6734 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6735 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6736 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6737 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6738 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6739 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6740 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6741 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6742 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6743 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6744 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6745 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6746 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6747 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6748 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6749 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6750 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6751 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6752 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6753 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6754 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6755 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6756 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6757 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6758 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6759 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6760 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6761 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6762 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6763 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6764 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6765 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6766 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6767 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6768 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6769 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6770 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6771 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6772 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6773 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6774 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6775 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6776 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6777 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6778 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6779 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6780 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6781 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6782 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6783 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6784 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6785 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6786 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6787 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6788 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6789 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6790 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6791 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6792 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6793 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6794 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6795 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6796 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6797 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6798 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6799 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6800 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6801 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6802 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6803 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6804 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6805 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6806 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6807 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6808 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6809 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6810 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6811 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6812 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6813 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6814 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6815 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6816 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6817 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6818 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6819 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6820 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6821 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6822 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6823 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6824 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6825 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6826 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6827 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6828 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6829 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6830 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6831 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6832 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6833 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6834 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6835 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6836 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6837 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6838 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6839 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6840 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6841 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6842 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6843 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6844 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6845 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6846 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6847 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6848 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6849 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6850 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6851 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6852 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6853 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6854 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6855 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6856 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6857 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6858 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6859 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6860 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6861 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6862 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6863 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6864 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6865 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6866 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6867 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6868 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6869 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6870 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6871 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6872 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6873 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6874 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6875 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6876 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6877 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6878 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6879 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6880 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6881 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6882 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6883 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6884 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6885 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6886 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6887 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6888 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6889 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6890 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6891 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6892 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6893 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6894 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6895 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6896 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6897 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6898 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6899 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6900 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6901 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6902 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6903 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6904 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6905 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6906 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6907 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6908 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6909 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6910 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6911 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6912 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6913 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6914 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6915 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6916 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6917 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6918 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6919 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6920 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6921 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6922 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6923 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6924 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6925 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6926 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6927 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6928 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6929 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6930 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6931 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6932 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6933 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6934 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6935 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6936 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6937 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6938 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6939 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6940 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6941 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6942 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6943 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6944 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6945 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6946 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6947 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6948 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6949 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6950 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6951 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6952 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6953 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6954 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6955 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6956 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6957 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6958 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6959 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6960 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6961 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6962 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6963 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6964 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6965 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6966 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6967 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6968 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6969 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6970 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6971 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6972 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6973 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6974 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6975 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6976 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6977 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6978 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6979 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6980 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6981 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6982 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6983 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6984 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6985 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6986 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6987 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6988 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6989 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6990 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6991 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6992 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6993 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6994 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6995 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6996 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6997 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6998 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		6999 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7000 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7001 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7002 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7003 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7004 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7005 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7006 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7007 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7008 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7009 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7010 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7011 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7012 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7013 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7014 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7015 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7016 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7017 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7018 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7019 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7020 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7021 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7022 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7023 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7024 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7025 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7026 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7027 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7028 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7029 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7030 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7031 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7032 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7033 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7034 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7035 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7036 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7037 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7038 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7039 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7040 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7041 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7042 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7043 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7044 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7045 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7046 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7047 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7048 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7049 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7050 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7051 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7052 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7053 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7054 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7055 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7056 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7057 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7058 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7059 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7060 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7061 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7062 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7063 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7064 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7065 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7066 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7067 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7068 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7069 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7070 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7071 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7072 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7073 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7074 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7075 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7076 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7077 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7078 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7079 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7080 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7081 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7082 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7083 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7084 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7085 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7086 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7087 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7088 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7089 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7090 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7091 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7092 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7093 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7094 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7095 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7096 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7097 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7098 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7099 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7100 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7101 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7102 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7103 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7104 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7105 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7106 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7107 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7108 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7109 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7110 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7111 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7112 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7113 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7114 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7115 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7116 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7117 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7118 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7119 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7120 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7121 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7122 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7123 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7124 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7125 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7126 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7127 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7128 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7129 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7130 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7131 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7132 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7133 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7134 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7135 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7136 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7137 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7138 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7139 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7140 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7141 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7142 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7143 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7144 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7145 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7146 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7147 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7148 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7149 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7150 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7151 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7152 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7153 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7154 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7155 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7156 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7157 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7158 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7159 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7160 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7161 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7162 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7163 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7164 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7165 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7166 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7167 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7168 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7169 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7170 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7171 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7172 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7173 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7174 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7175 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7176 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7177 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7178 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7179 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7180 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7181 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7182 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7183 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7184 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7185 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7186 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7187 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7188 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7189 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7190 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7191 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7192 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7193 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7194 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7195 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7196 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7197 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7198 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7199 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7200 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7201 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7202 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7203 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7204 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7205 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7206 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7207 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7208 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7209 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7210 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7211 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7212 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7213 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7214 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7215 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7216 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7217 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7218 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7219 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7220 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7221 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7222 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7223 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7224 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7225 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7226 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7227 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7228 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7229 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7230 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7231 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7232 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7233 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7234 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7235 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7236 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7237 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7238 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7239 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7240 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7241 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7242 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7243 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7244 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7245 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7246 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7247 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7248 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7249 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7250 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7251 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7252 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7253 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7254 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7255 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7256 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7257 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7258 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7259 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7260 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7261 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7262 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7263 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7264 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7265 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7266 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7267 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7268 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7269 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7270 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7271 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7272 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7273 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7274 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7275 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7276 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7277 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7278 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7279 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7280 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7281 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7282 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7283 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7284 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7285 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7286 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7287 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7288 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7289 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7290 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7291 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7292 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7293 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7294 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7295 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7296 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7297 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7298 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7299 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7300 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7301 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7302 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7303 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7304 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7305 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7306 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7307 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7308 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7309 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7310 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7311 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7312 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7313 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7314 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7315 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7316 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7317 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7318 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7319 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7320 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7321 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7322 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7323 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7324 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7325 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7326 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7327 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7328 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7329 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7330 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7331 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7332 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7333 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7334 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7335 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7336 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7337 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7338 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7339 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7340 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7341 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7342 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7343 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7344 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7345 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7346 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7347 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7348 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7349 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7350 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7351 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7352 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7353 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7354 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7355 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7356 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7357 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7358 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7359 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7360 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7361 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7362 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7363 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7364 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7365 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7366 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7367 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7368 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7369 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7370 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7371 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7372 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7373 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7374 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7375 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7377 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7378 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7379 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7380 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7381 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7382 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7383 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7384 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7385 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7386 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7387 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7388 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7389 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7390 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7391 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7392 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7393 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7394 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7395 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7396 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7397 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7398 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7399 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7400 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7401 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7402 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7403 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7404 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7405 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7406 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7407 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7408 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7409 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7410 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7411 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7412 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7413 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7414 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7415 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7416 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7417 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7418 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7419 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7420 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7421 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7422 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7423 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7424 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7425 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7426 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7427 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7428 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7429 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7430 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7431 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7432 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7433 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7434 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7435 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7436 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7437 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7438 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7439 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7440 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7441 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7442 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7443 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7444 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7445 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7446 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7447 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7448 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7449 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7450 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7451 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7452 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7453 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7454 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7455 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7456 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7457 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7458 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7459 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7460 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7461 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7462 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7463 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7464 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7465 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7466 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7467 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7468 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7469 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7470 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7471 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7472 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7473 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7474 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7475 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7476 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7477 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7478 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7479 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7480 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7481 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7482 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7483 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7484 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7485 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7486 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7487 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7488 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7489 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7490 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7491 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7492 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7493 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7494 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7495 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7496 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7497 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7498 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7499 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7500 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7501 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7502 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7503 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7504 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7505 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7506 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7507 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7508 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7509 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7510 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7511 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7512 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7513 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7514 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7515 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7516 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7517 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7518 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7519 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7520 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7521 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7522 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7523 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7524 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7525 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7526 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7527 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7528 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7529 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7530 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7531 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7532 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7533 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7534 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7535 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7536 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7537 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7538 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7539 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7540 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7541 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7542 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7543 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7544 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7545 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7546 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7547 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7548 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7549 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7550 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7551 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7552 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7553 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7554 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7555 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7556 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7557 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7558 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7559 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7560 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7561 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7562 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7563 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7564 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7565 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7566 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7567 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7568 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7569 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7570 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7571 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7572 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7573 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7574 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7575 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7576 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7577 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7578 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7579 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7580 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7581 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7582 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7583 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7584 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7585 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7586 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7587 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7588 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7589 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7590 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7591 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7592 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7593 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7594 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7595 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7596 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7597 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7598 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7599 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7600 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7601 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7602 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7603 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7604 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7605 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7606 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7607 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7608 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7609 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7610 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7611 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7612 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7613 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7614 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7615 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7616 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7617 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7618 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7619 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7620 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7621 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7622 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7623 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7624 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7625 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7626 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7627 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7628 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7629 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7630 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7631 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7632 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7633 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7634 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7635 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7636 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7637 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7638 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7639 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7640 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7641 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7642 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7643 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7644 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7645 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7646 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7647 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7648 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7649 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7650 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7651 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7652 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7653 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7654 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7655 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7656 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7657 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7658 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7659 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7660 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7661 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7662 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7663 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7664 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7665 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7666 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7667 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7668 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7669 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7670 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7671 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7672 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7673 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7674 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7675 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7676 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7677 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7678 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7679 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7680 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7681 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7682 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7683 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7684 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7685 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7686 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7687 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7688 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7689 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7690 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7691 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7692 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7693 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7694 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7695 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7696 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7697 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7698 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7699 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7700 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7701 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7702 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7703 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7704 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7705 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7706 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7707 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7708 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7709 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7710 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7711 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7712 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7713 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7714 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7715 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7716 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7717 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7718 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7719 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7720 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7721 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7722 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7723 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7724 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7725 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7726 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7727 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7728 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7729 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7730 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7731 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7732 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7733 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7734 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7735 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7736 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7737 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7738 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7739 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7740 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7741 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7742 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7743 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7744 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7745 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7746 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7747 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7748 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7749 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7750 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7751 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7752 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7753 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7754 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7755 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7756 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7757 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7758 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7759 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7760 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7761 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7762 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7763 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7764 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7765 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7766 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7767 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7768 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7769 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7770 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7771 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7772 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7773 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7774 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7775 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7776 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7777 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7778 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7779 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7780 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7781 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7782 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7783 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7784 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7785 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7786 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7787 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7788 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7789 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7790 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7791 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7792 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7793 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7794 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7795 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7796 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7797 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7798 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7799 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7800 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7801 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7802 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7803 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7804 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7805 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7806 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7807 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7808 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7809 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7810 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7811 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7812 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7813 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7814 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7815 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7816 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7817 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7818 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7819 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7820 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7821 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7822 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7823 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7824 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7825 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7826 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7827 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7828 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7829 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7830 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7831 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7832 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7833 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7834 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7835 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7836 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7837 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7838 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7839 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7840 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7841 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7842 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7843 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7844 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7845 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7846 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7847 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7848 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7849 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7850 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7851 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7852 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7853 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7854 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7855 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7856 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7857 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7858 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7859 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7860 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7861 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7862 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7863 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7864 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7865 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7866 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7867 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7868 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7869 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7870 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7871 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7872 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7873 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7874 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7875 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7876 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7877 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7878 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7879 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7880 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7881 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7882 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7883 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7884 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7885 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7886 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7887 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7888 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7889 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7890 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7891 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7892 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7893 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7894 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7895 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7896 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7897 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7898 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7899 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7900 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7901 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7902 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7903 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7904 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7905 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7906 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7907 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7908 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7909 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7910 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7911 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7912 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7913 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7914 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7915 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7916 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7917 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7918 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7919 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7920 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7921 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7922 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7923 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7924 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7925 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7926 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7927 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7928 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7929 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7930 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7931 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7932 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7933 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7934 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7935 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7936 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7937 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7938 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7939 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7940 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7941 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7942 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7943 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7944 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7945 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7946 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7947 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7948 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7949 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7950 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7951 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7952 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7953 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7954 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7955 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7956 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7957 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7958 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7959 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7960 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7961 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7962 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7963 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7964 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7965 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7966 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7967 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7968 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7969 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7970 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7971 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7972 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7973 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7974 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7975 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7976 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7977 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7978 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7979 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7980 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7981 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7982 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7983 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7984 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7985 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7986 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7987 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7988 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7989 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7990 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7991 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7992 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7993 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7994 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7995 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7996 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7997 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7998 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		7999 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8000 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8001 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8002 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8003 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8004 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8005 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8006 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8007 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8008 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8009 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8010 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8011 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8012 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8013 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8014 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8015 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8016 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8017 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8018 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8019 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8020 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8021 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8022 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8023 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8024 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8025 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8026 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8027 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8028 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8029 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8030 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8031 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8032 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8033 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8034 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8035 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8036 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8037 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8038 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8039 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8040 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8041 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8042 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8043 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8044 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8045 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8046 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8047 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8048 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8049 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8050 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8051 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8052 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8053 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8054 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8055 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8056 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8057 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8058 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8059 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8060 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8061 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8062 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8063 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8064 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8065 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8066 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8067 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8068 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8069 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8070 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8071 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8072 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8073 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8074 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8075 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8076 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8077 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8078 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8079 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8080 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8081 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8082 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8083 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8084 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8085 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8086 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8087 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8088 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8089 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8090 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8091 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8092 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8093 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8094 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8095 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8096 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8097 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8098 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8099 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8100 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8101 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8102 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8103 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8104 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8105 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8106 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8107 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8108 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8109 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8110 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8111 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8112 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8113 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8114 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8115 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8116 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8117 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8118 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8119 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8120 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8121 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8122 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8123 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8124 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8125 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8126 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8127 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8128 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8129 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8130 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8131 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8132 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8133 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8134 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8135 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8136 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8137 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8138 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8139 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8140 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8141 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8142 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8143 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8144 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8145 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8146 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8147 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8148 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8149 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8150 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8151 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8152 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8153 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8154 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8155 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8156 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8157 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8158 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8159 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8160 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8161 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8162 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8163 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8164 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8165 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8166 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8167 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8168 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8169 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8170 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8171 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8172 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8173 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8174 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8175 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8176 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8177 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8178 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8179 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8180 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8181 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8182 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8183 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8184 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8185 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8186 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8187 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8188 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8189 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8190 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8191 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8192 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8193 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8194 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8195 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8196 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8197 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8198 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8199 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8200 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8201 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8202 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8203 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8204 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8205 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8206 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8207 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8208 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8209 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8210 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8211 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8212 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8213 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8214 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8215 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8216 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8217 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8218 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8219 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8220 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8221 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8222 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8223 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8224 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8225 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8226 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8227 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8228 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8229 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8230 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8231 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8232 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8233 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8234 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8235 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8236 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8237 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8238 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8239 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8240 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8241 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8242 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8243 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8244 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8245 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8246 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8247 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8248 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8249 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8250 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8251 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8252 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8253 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8254 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8255 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8256 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8257 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8258 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8259 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8260 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8261 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8262 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8263 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8264 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8265 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8266 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8267 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8268 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8269 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8270 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8271 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8272 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8273 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8274 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8275 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8276 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8277 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8278 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8279 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8280 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8281 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8282 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8283 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8284 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8285 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8286 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8287 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8288 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8289 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8290 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8291 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8292 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8293 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8294 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8295 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8296 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8297 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8298 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8299 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8300 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8301 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8302 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8303 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8304 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8305 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8306 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8307 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8308 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8309 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8310 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8311 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8312 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8313 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8314 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8315 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8316 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8317 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8318 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8319 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8320 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8321 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8322 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8323 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8324 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8325 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8326 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8327 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8328 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8329 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8330 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8331 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8332 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8333 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8334 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8335 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8336 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8337 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8338 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8339 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8340 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8341 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8342 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8343 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8344 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8345 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8346 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8347 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8348 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8349 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8350 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8351 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8352 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8353 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8354 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8355 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8356 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8357 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8358 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8359 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8360 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8361 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8362 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8363 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8364 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8365 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8366 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8367 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8368 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8369 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8370 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8371 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8372 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8373 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8374 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8375 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8377 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8378 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8379 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8380 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8381 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8382 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8383 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8384 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8385 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8386 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8387 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8388 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8389 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8390 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8391 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8392 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8393 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8394 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8395 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8396 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8397 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8398 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8399 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8400 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8401 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8402 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8403 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8404 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8405 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8406 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8407 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8408 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8409 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8410 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8411 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8412 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8413 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8414 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8415 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8416 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8417 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8418 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8419 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8420 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8421 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8422 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8423 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8424 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8425 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8426 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8427 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8428 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8429 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8430 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8431 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8432 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8433 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8434 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8435 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8436 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8437 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8438 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8439 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8440 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8441 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8442 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8443 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8444 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8445 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8446 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8447 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8448 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8449 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8450 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8451 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8452 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8453 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8454 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8455 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8456 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8457 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8458 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8459 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8460 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8461 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8462 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8463 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8464 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8465 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8466 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8467 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8468 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8469 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8470 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8471 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8472 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8473 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8474 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8475 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8476 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8477 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8478 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8479 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8480 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8481 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8482 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8483 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8484 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8485 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8486 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8487 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8488 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8489 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8490 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8491 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8492 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8493 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8494 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8495 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8496 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8497 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8498 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8499 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8500 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8501 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8502 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8503 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8504 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8505 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8506 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8507 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8508 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8509 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8510 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8511 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8512 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8513 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8514 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8515 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8516 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8517 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8518 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8519 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8520 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8521 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8522 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8523 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8524 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8525 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8526 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8527 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8528 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8529 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8530 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8531 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8532 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8533 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8534 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8535 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8536 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8537 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8538 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8539 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8540 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8541 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8542 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8543 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8544 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8545 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8546 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8547 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8548 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8549 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8550 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8551 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8552 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8553 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8554 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8555 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8556 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8557 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8558 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8559 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8560 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8561 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8562 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8563 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8564 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8565 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8566 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8567 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8568 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8569 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8570 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8571 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8572 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8573 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8574 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8575 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8576 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8577 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8578 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8579 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8580 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8581 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8582 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8583 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8584 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8585 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8586 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8587 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8588 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8589 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8590 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8591 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8592 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8593 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8594 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8595 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8596 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8597 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8598 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8599 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8600 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8601 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8602 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8603 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8604 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8605 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8606 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8607 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8608 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8609 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8610 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8611 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8612 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8613 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8614 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8615 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8616 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8617 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8618 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8619 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8620 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8621 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8622 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8623 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8624 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8625 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8626 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8627 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8628 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8629 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8630 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8631 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8632 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8633 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8634 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8635 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8636 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8637 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8638 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8639 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8640 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8641 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8642 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8643 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8644 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8645 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8646 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8647 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8648 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8649 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8650 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8651 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8652 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8653 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8654 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8655 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8656 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8657 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8658 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8659 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8660 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8661 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8662 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8663 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8664 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8665 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8666 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8667 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8668 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8669 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8670 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8671 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8672 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8673 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8674 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8675 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8676 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8677 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8678 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8679 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8680 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8681 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8682 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8683 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8684 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8685 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8686 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8687 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8688 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8689 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8690 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8691 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8692 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8693 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8694 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8695 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8696 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8697 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8698 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8699 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8700 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8701 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8702 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8703 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8704 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8705 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8706 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8707 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8708 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8709 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8710 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8711 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8712 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8713 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8714 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8715 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8716 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8717 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8718 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8719 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8720 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8721 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8722 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8723 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8724 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8725 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8726 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8727 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8728 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8729 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8730 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8731 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8732 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8733 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8734 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8735 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8736 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8737 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8738 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8739 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8740 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8741 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8742 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8743 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8744 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8745 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8746 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8747 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8748 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8749 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8750 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8751 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8752 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8753 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8754 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8755 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8756 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8757 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8758 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8759 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8760 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8761 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8762 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8763 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8764 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8765 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8766 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8767 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8768 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8769 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8770 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8771 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8772 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8773 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8774 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8775 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8776 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8777 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8778 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8779 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8780 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8781 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8782 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8783 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8784 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8785 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8786 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8787 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8788 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8789 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8790 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8791 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8792 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8793 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8794 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8795 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8796 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8797 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8798 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8799 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8800 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8801 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8802 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8803 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8804 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8805 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8806 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8807 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8808 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8809 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8810 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8811 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8812 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8813 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8814 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8815 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8816 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8817 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8818 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8819 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8820 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8821 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8822 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8823 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8824 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8825 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8826 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8827 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8828 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8829 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8830 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8831 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8832 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8833 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8834 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8835 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8836 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8837 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8838 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8839 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8840 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8841 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8842 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8843 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8844 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8845 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8846 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8847 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8848 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8849 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8850 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8851 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8852 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8853 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8854 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8855 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8856 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8857 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8858 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8859 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8860 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8861 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8862 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8863 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8864 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8865 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8866 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8867 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8868 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8869 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8870 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8871 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8872 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8873 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8874 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8875 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8876 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8877 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8878 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8879 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8880 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8881 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8882 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8883 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8884 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8885 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8886 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8887 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8888 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8889 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8890 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8891 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8892 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8893 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8894 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8895 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8896 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8897 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8898 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8899 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8900 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8901 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8902 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8903 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8904 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8905 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8906 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8907 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8908 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8909 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8910 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8911 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8912 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8913 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8914 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8915 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8916 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8917 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8918 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8919 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8920 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8921 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8922 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8923 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8924 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8925 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8926 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8927 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8928 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8929 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8930 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8931 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8932 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8933 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8934 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8935 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8936 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8937 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8938 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8939 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8940 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8941 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8942 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8943 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8944 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8945 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8946 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8947 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8948 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8949 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8950 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8951 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8952 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8953 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8954 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8955 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8956 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8957 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8958 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8959 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8960 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8961 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8962 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8963 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8964 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8965 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8966 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8967 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8968 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8969 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8970 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8971 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8972 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8973 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8974 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8975 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8976 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8977 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8978 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8979 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8980 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8981 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8982 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8983 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8984 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8985 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8986 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8987 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8988 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8989 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8990 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8991 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8992 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8993 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8994 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8995 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8996 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8997 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8998 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		8999 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9000 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9001 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9002 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9003 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9004 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9005 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9006 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9007 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9008 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9009 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9010 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9011 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9012 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9013 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9014 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9015 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9016 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9017 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9018 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9019 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9020 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9021 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9022 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9023 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9024 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9025 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9026 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9027 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9028 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9029 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9030 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9031 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9032 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9033 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9034 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9035 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9036 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9037 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9038 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9039 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9040 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9041 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9042 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9043 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9044 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9045 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9046 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9047 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9048 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9049 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9050 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9051 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9052 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9053 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9054 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9055 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9056 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9057 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9058 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9059 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9060 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9061 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9062 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9063 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9064 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9065 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9066 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9067 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9068 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9069 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9070 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9071 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9072 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9073 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9074 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9075 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9076 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9077 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9078 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9079 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9080 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9081 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9082 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9083 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9084 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9085 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9086 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9087 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9088 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9089 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9090 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9091 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9092 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9093 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9094 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9095 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9096 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9097 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9098 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9099 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9100 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9101 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9102 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9103 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9104 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9105 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9106 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9107 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9108 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9109 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9110 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9111 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9112 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9113 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9114 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9115 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9116 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9117 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9118 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9119 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9120 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9121 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9122 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9123 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9124 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9125 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9126 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9127 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9128 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9129 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9130 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9131 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9132 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9133 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9134 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9135 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9136 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9137 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9138 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9139 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9140 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9141 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9142 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9143 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9144 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9145 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9146 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9147 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9148 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9149 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9150 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9151 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9152 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9153 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9154 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9155 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9156 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9157 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9158 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9159 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9160 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9161 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9162 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9163 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9164 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9165 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9166 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9167 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9168 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9169 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9170 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9171 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9172 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9173 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9174 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9175 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9176 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9177 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9178 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9179 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9180 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9181 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9182 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9183 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9184 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9185 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9186 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9187 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9188 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9189 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9190 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9191 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9192 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9193 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9194 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9195 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9196 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9197 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9198 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9199 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9200 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9201 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9202 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9203 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9204 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9205 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9206 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9207 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9208 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9209 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9210 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9211 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9212 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9213 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9214 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9215 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9216 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9217 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9218 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9219 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9220 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9221 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9222 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9223 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9224 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9225 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9226 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9227 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9228 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9229 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9230 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9231 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9232 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9233 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9234 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9235 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9236 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9237 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9238 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9239 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9240 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9241 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9242 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9243 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9244 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9245 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9246 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9247 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9248 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9249 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9250 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9251 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9252 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9253 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9254 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9255 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9256 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9257 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9258 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9259 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9260 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9261 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9262 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9263 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9264 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9265 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9266 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9267 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9268 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9269 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9270 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9271 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9272 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9273 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9274 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9275 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9276 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9277 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9278 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9279 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9280 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9281 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9282 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9283 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9284 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9285 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9286 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9287 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9288 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9289 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9290 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9291 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9292 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9293 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9294 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9295 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9296 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9297 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9298 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9299 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9300 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9301 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9302 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9303 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9304 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9305 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9306 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9307 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9308 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9309 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9310 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9311 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9312 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9313 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9314 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9315 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9316 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9317 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9318 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9319 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9320 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9321 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9322 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9323 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9324 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9325 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9326 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9327 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9328 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9329 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9330 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9331 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9332 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9333 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9334 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9335 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9336 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9337 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9338 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9339 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9340 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9341 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9342 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9343 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9344 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9345 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9346 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9347 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9348 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9349 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9350 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9351 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9352 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9353 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9354 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9355 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9356 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9357 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9358 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9359 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9360 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9361 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9362 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9363 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9364 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9365 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9366 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9367 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9368 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9369 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9370 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9371 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9372 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9373 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9374 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9375 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9377 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9378 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9379 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9380 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9381 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9382 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9383 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9384 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9385 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9386 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9387 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9388 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9389 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9390 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9391 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9392 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9393 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9394 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9395 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9396 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9397 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9398 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9399 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9400 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9401 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9402 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9403 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9404 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9405 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9406 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9407 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9408 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9409 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9410 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9411 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9412 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9413 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9414 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9415 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9416 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9417 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9418 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9419 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9420 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9421 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9422 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9423 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9424 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9425 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9426 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9427 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9428 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9429 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9430 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9431 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9432 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9433 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9434 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9435 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9436 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9437 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9438 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9439 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9440 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9441 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9442 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9443 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9444 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9445 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9446 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9447 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9448 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9449 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9450 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9451 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9452 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9453 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9454 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9455 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9456 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9457 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9458 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9459 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9460 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9461 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9462 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9463 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9464 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9465 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9466 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9467 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9468 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9469 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9470 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9471 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9472 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9473 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9474 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9475 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9476 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9477 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9478 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9479 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9480 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9481 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9482 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9483 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9484 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9485 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9486 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9487 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9488 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9489 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9490 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9491 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9492 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9493 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9494 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9495 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9496 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9497 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9498 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9499 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9500 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9501 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9502 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9503 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9504 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9505 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9506 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9507 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9508 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9509 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9510 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9511 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9512 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9513 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9514 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9515 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9516 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9517 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9518 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9519 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9520 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9521 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9522 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9523 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9524 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9525 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9526 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9527 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9528 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9529 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9530 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9531 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9532 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9533 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9534 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9535 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9536 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9537 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9538 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9539 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9540 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9541 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9542 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9543 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9544 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9545 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9546 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9547 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9548 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9549 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9550 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9551 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9552 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9553 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9554 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9555 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9556 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9557 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9558 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9559 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9560 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9561 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9562 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9563 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9564 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9565 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9566 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9567 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9568 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9569 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9570 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9571 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9572 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9573 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9574 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9575 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9576 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9577 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9578 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9579 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9580 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9581 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9582 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9583 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9584 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9585 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9586 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9587 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9588 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9589 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9590 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9591 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9592 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9593 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9594 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9595 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9596 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9597 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9598 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9599 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9600 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9601 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9602 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9603 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9604 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9605 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9606 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9607 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9608 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9609 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9610 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9611 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9612 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9613 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9614 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9615 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9616 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9617 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9618 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9619 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9620 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9621 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9622 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9623 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9624 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9625 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9626 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9627 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9628 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9629 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9630 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9631 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9632 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9633 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9634 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9635 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9636 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9637 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9638 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9639 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9640 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9641 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9642 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9643 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9644 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9645 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9646 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9647 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9648 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9649 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9650 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9651 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9652 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9653 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9654 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9655 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9656 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9657 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9658 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9659 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9660 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9661 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9662 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9663 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9664 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9665 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9666 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9667 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9668 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9669 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9670 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9671 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9672 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9673 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9674 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9675 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9676 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9677 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9678 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9679 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9680 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9681 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9682 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9683 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9684 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9685 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9686 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9687 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9688 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9689 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9690 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9691 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9692 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9693 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9694 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9695 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9696 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9697 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9698 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9699 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9700 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9701 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9702 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9703 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9704 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9705 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9706 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9707 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9708 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9709 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9710 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9711 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9712 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9713 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9714 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9715 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9716 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9717 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9718 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9719 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9720 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9721 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9722 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9723 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9724 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9725 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9726 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9727 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9728 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9729 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9730 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9731 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9732 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9733 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9734 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9735 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9736 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9737 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9738 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9739 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9740 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9741 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9742 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9743 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9744 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9745 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9746 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9747 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9748 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9749 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9750 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9751 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9752 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9753 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9754 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9755 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9756 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9757 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9758 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9759 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9760 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9761 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9762 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9763 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9764 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9765 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9766 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9767 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9768 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9769 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9770 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9771 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9772 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9773 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9774 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9775 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9776 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9777 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9778 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9779 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9780 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9781 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9782 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9783 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9784 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9785 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9786 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9787 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9788 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9789 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9790 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9791 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9792 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9793 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9794 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9795 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9796 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9797 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9798 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9799 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9800 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9801 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9802 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9803 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9804 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9805 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9806 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9807 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9808 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9809 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9810 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9811 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9812 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9813 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9814 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9815 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9816 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9817 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9818 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9819 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9820 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9821 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9822 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9823 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9824 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9825 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9826 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9827 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9828 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9829 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9830 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9831 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9832 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9833 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9834 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9835 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9836 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9837 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9838 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9839 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9840 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9841 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9842 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9843 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9844 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9845 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9846 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9847 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9848 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9849 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9850 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9851 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9852 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9853 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9854 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9855 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9856 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9857 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9858 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9859 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9860 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9861 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9862 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9863 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9864 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9865 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9866 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9867 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9868 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9869 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9870 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9871 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9872 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9873 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9874 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9875 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9876 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9877 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9878 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9879 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9880 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9881 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9882 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9883 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9884 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9885 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9886 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9887 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9888 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9889 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9890 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9891 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9892 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9893 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9894 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9895 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9896 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9897 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9898 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9899 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9900 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9901 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9902 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9903 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9904 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9905 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9906 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9907 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9908 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9909 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9910 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9911 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9912 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9913 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9914 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9915 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9916 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9917 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9918 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9919 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9920 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9921 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9922 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9923 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9924 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9925 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9926 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9927 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9928 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9929 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9930 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9931 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9932 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9933 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9934 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9935 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9936 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9937 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9938 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9939 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9940 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9941 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9942 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9943 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9944 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9945 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9946 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9947 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9948 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9949 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9950 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9951 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9952 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9953 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9954 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9955 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9956 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9957 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9958 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9959 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9960 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9961 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9962 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9963 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9964 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9965 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9966 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9967 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9968 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9969 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9970 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9971 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9972 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9973 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9974 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9975 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9976 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9977 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9978 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9979 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9980 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9981 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9982 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9983 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9984 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9985 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9986 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9987 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9988 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9989 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9990 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9991 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9992 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9993 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9994 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9995 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9996 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9997 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9998 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		9999 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10000 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10001 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10002 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10003 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10004 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10005 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10006 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10007 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10008 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10009 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10010 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10011 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10012 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10013 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10014 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10015 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10016 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10017 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10018 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10019 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10020 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10021 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10022 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10023 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10024 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10025 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10026 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10027 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10028 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10029 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10030 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10031 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10032 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10033 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10034 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10035 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10036 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10037 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10038 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10039 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10040 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10041 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10042 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10043 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10044 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10045 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10046 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10047 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10048 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10049 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10050 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10051 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10052 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10053 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10054 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10055 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10056 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10057 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10058 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10059 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10060 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10061 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10062 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10063 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10064 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10065 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10066 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10067 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10068 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10069 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10070 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10071 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10072 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10073 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10074 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10075 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10076 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10077 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10078 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10079 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10080 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10081 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10082 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10083 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10084 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10085 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10086 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10087 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10088 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10089 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10090 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10091 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10092 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10093 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10094 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10095 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10096 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10097 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10098 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10099 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10100 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10101 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10102 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10103 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10104 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10105 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10106 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10107 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10108 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10109 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10110 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10111 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10112 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10113 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10114 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10115 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10116 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10117 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10118 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10119 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10120 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10121 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10122 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10123 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10124 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10125 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10126 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10127 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10128 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10129 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10130 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10131 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10132 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10133 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10134 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10135 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10136 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10137 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10138 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10139 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10140 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10141 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10142 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10143 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10144 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10145 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10146 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10147 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10148 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10149 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10150 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10151 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10152 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10153 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10154 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10155 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10156 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10157 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10158 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10159 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10160 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10161 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10162 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10163 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10164 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10165 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10166 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10167 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10168 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10169 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10170 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10171 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10172 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10173 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10174 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10175 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10176 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10177 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10178 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10179 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10180 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10181 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10182 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10183 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10184 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10185 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10186 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10187 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10188 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10189 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10190 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10191 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10192 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10193 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10194 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10195 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10196 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10197 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10198 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10199 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10200 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10201 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10202 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10203 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10204 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10205 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10206 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10207 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10208 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10209 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10210 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10211 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10212 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10213 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10214 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10215 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10216 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10217 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10218 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10219 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10220 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10221 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10222 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10223 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10224 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10225 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10226 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10227 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10228 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10229 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10230 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10231 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10232 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10233 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10234 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10235 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10236 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10237 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10238 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10239 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10240 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10241 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10242 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10243 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10244 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10245 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10246 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10247 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10248 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10249 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10250 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10251 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10252 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10253 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10254 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10255 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10256 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10257 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10258 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10259 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10260 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10261 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10262 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10263 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10264 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10265 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10266 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10267 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10268 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10269 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10270 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10271 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10272 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10273 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10274 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10275 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10276 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10277 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10278 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10279 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10280 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10281 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10282 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10283 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10284 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10285 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10286 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10287 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10288 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10289 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10290 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10291 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10292 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10293 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10294 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10295 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10296 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10297 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10298 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10299 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10300 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10301 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10302 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		10303 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		others => x"00000000"
	);

begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;