
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER
-- DATE: Thu May 31 11:44:22 2018

	signal mem : ram_t := (
	
--			***** COLOR PALLETE *****

		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00277FFF", -- R: 255 G: 127 B: 39
		2 =>	x"004798FF", -- R: 255 G: 152 B: 71
		3 =>	x"000000FF", -- R: 255 G: 0 B: 0
		4 =>	x"007F7F7F", -- R: 127 G: 127 B: 127
		5 =>	x"00FF0000", -- R: 0 G: 0 B: 255
		6 =>	x"0000FFFF", -- R: 255 G: 255 B: 0
		7 =>	x"00007F00", -- R: 0 G: 127 B: 0
		8 =>	x"004C4C4C", -- R: 76 G: 76 B: 76
		9 =>	x"007F007F", -- R: 127 G: 0 B: 127
		10 =>	x"0000007F", -- R: 127 G: 0 B: 0
		11 =>	x"00007F82", -- R: 130 G: 127 B: 0
		12 =>	x"00666666", -- R: 102 G: 102 B: 102
		13 =>	x"009800FF", -- R: 255 G: 0 B: 152
		14 =>	x"009800A4", -- R: 164 G: 0 B: 152
		15 =>	x"00980000", -- R: 0 G: 0 B: 152
		16 =>	x"005480D7", -- R: 215 G: 128 B: 84
		17 =>	x"00862138", -- R: 56 G: 33 B: 134
		18 =>	x"00990000", -- R: 0 G: 0 B: 153
		19 =>	x"00862136", -- R: 54 G: 33 B: 134
		20 =>	x"00980124", -- R: 36 G: 1 B: 152
		21 =>	x"00980095", -- R: 149 G: 0 B: 152
		22 =>	x"009800A5", -- R: 165 G: 0 B: 152
		23 =>	x"00980094", -- R: 148 G: 0 B: 152
		24 =>	x"009800DF", -- R: 223 G: 0 B: 152
		25 =>	x"009800A7", -- R: 167 G: 0 B: 152
		26 =>	x"0098016B", -- R: 107 G: 1 B: 152
		27 =>	x"00000000", -- Unused
		28 =>	x"00000000", -- Unused
		29 =>	x"00000000", -- Unused
		30 =>	x"00000000", -- Unused
		31 =>	x"00000000", -- Unused
		32 =>	x"00000000", -- Unused
		33 =>	x"00000000", -- Unused
		34 =>	x"00000000", -- Unused
		35 =>	x"00000000", -- Unused
		36 =>	x"00000000", -- Unused
		37 =>	x"00000000", -- Unused
		38 =>	x"00000000", -- Unused
		39 =>	x"00000000", -- Unused
		40 =>	x"00000000", -- Unused
		41 =>	x"00000000", -- Unused
		42 =>	x"00000000", -- Unused
		43 =>	x"00000000", -- Unused
		44 =>	x"00000000", -- Unused
		45 =>	x"00000000", -- Unused
		46 =>	x"00000000", -- Unused
		47 =>	x"00000000", -- Unused
		48 =>	x"00000000", -- Unused
		49 =>	x"00000000", -- Unused
		50 =>	x"00000000", -- Unused
		51 =>	x"00000000", -- Unused
		52 =>	x"00000000", -- Unused
		53 =>	x"00000000", -- Unused
		54 =>	x"00000000", -- Unused
		55 =>	x"00000000", -- Unused
		56 =>	x"00000000", -- Unused
		57 =>	x"00000000", -- Unused
		58 =>	x"00000000", -- Unused
		59 =>	x"00000000", -- Unused
		60 =>	x"00000000", -- Unused
		61 =>	x"00000000", -- Unused
		62 =>	x"00000000", -- Unused
		63 =>	x"00000000", -- Unused
		64 =>	x"00000000", -- Unused
		65 =>	x"00000000", -- Unused
		66 =>	x"00000000", -- Unused
		67 =>	x"00000000", -- Unused
		68 =>	x"00000000", -- Unused
		69 =>	x"00000000", -- Unused
		70 =>	x"00000000", -- Unused
		71 =>	x"00000000", -- Unused
		72 =>	x"00000000", -- Unused
		73 =>	x"00000000", -- Unused
		74 =>	x"00000000", -- Unused
		75 =>	x"00000000", -- Unused
		76 =>	x"00000000", -- Unused
		77 =>	x"00000000", -- Unused
		78 =>	x"00000000", -- Unused
		79 =>	x"00000000", -- Unused
		80 =>	x"00000000", -- Unused
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
		255 =>	x"00000000", -- Unused

--			***** 16x16 IMAGES *****


		256 =>	x"01010101", -- IMG_16x16_background
		257 =>	x"01010101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01010101",
		261 =>	x"01010101",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01010101",
		265 =>	x"01010101",
		266 =>	x"01010101",
		267 =>	x"01010101",
		268 =>	x"01010101",
		269 =>	x"01010101",
		270 =>	x"01010101",
		271 =>	x"01010101",
		272 =>	x"01010101",
		273 =>	x"01010101",
		274 =>	x"01010101",
		275 =>	x"01010101",
		276 =>	x"01010101",
		277 =>	x"01010101",
		278 =>	x"01010101",
		279 =>	x"01010101",
		280 =>	x"01010101",
		281 =>	x"01010101",
		282 =>	x"01010101",
		283 =>	x"01010101",
		284 =>	x"01010101",
		285 =>	x"01010101",
		286 =>	x"01010101",
		287 =>	x"01010101",
		288 =>	x"01010101",
		289 =>	x"01010101",
		290 =>	x"01010101",
		291 =>	x"01010101",
		292 =>	x"01010101",
		293 =>	x"01010101",
		294 =>	x"01010101",
		295 =>	x"01010101",
		296 =>	x"01010101",
		297 =>	x"01010101",
		298 =>	x"01010101",
		299 =>	x"01010101",
		300 =>	x"01010101",
		301 =>	x"01010101",
		302 =>	x"01010101",
		303 =>	x"01010101",
		304 =>	x"01010101",
		305 =>	x"01010101",
		306 =>	x"01010101",
		307 =>	x"01010101",
		308 =>	x"01010101",
		309 =>	x"01010101",
		310 =>	x"01010101",
		311 =>	x"01010101",
		312 =>	x"01010101",
		313 =>	x"01010101",
		314 =>	x"01010101",
		315 =>	x"01010101",
		316 =>	x"01010101",
		317 =>	x"01010101",
		318 =>	x"01010101",
		319 =>	x"01010101",
		320 =>	x"02020202", -- IMG_16x16_bang
		321 =>	x"02020202",
		322 =>	x"02020302",
		323 =>	x"02020202",
		324 =>	x"02030302",
		325 =>	x"02020202",
		326 =>	x"02030303",
		327 =>	x"02030302",
		328 =>	x"02020303",
		329 =>	x"03030202",
		330 =>	x"03030303",
		331 =>	x"03030202",
		332 =>	x"02020303",
		333 =>	x"03030303",
		334 =>	x"03030303",
		335 =>	x"03030202",
		336 =>	x"00000003",
		337 =>	x"03000303",
		338 =>	x"00030300",
		339 =>	x"03000000",
		340 =>	x"00030003",
		341 =>	x"00030003",
		342 =>	x"00030300",
		343 =>	x"03000202",
		344 =>	x"00030003",
		345 =>	x"00030003",
		346 =>	x"00030300",
		347 =>	x"03000202",
		348 =>	x"00020003",
		349 =>	x"00030003",
		350 =>	x"00000300",
		351 =>	x"03000302",
		352 =>	x"00000303",
		353 =>	x"00000003",
		354 =>	x"00030000",
		355 =>	x"03000200",
		356 =>	x"00020003",
		357 =>	x"00030003",
		358 =>	x"00030300",
		359 =>	x"03000300",
		360 =>	x"00020003",
		361 =>	x"00030003",
		362 =>	x"00030300",
		363 =>	x"03000300",
		364 =>	x"00000003",
		365 =>	x"00030003",
		366 =>	x"00030300",
		367 =>	x"03000000",
		368 =>	x"02030303",
		369 =>	x"03020303",
		370 =>	x"03030303",
		371 =>	x"02020202",
		372 =>	x"02030303",
		373 =>	x"02020203",
		374 =>	x"03030302",
		375 =>	x"02020202",
		376 =>	x"03030202",
		377 =>	x"02020202",
		378 =>	x"03030202",
		379 =>	x"02020202",
		380 =>	x"02020202",
		381 =>	x"02020202",
		382 =>	x"03020202",
		383 =>	x"02020202",
		384 =>	x"00000000", -- IMG_16x16_car_blue
		385 =>	x"00000000",
		386 =>	x"00000000",
		387 =>	x"00000000",
		388 =>	x"00000404",
		389 =>	x"04000000",
		390 =>	x"00000000",
		391 =>	x"00000000",
		392 =>	x"00000404",
		393 =>	x"04000005",
		394 =>	x"00000000",
		395 =>	x"00000000",
		396 =>	x"00000004",
		397 =>	x"00000005",
		398 =>	x"05000000",
		399 =>	x"00000000",
		400 =>	x"00000505",
		401 =>	x"05050505",
		402 =>	x"05050000",
		403 =>	x"04040400",
		404 =>	x"00040405",
		405 =>	x"05050505",
		406 =>	x"05050505",
		407 =>	x"04040400",
		408 =>	x"00040404",
		409 =>	x"04060606",
		410 =>	x"05050505",
		411 =>	x"00040000",
		412 =>	x"00000505",
		413 =>	x"05060606",
		414 =>	x"06050505",
		415 =>	x"05050500",
		416 =>	x"00000505",
		417 =>	x"05060606",
		418 =>	x"06050505",
		419 =>	x"05050500",
		420 =>	x"00040404",
		421 =>	x"04060606",
		422 =>	x"05050505",
		423 =>	x"00040000",
		424 =>	x"00040405",
		425 =>	x"05050505",
		426 =>	x"05050505",
		427 =>	x"04040400",
		428 =>	x"00000505",
		429 =>	x"05050505",
		430 =>	x"05050000",
		431 =>	x"04040400",
		432 =>	x"00000004",
		433 =>	x"00000005",
		434 =>	x"05000000",
		435 =>	x"00000000",
		436 =>	x"00000404",
		437 =>	x"04000005",
		438 =>	x"00000000",
		439 =>	x"00000000",
		440 =>	x"00000404",
		441 =>	x"04000000",
		442 =>	x"00000000",
		443 =>	x"00000000",
		444 =>	x"00000000",
		445 =>	x"00000000",
		446 =>	x"00000000",
		447 =>	x"00000000",
		448 =>	x"02020202", -- IMG_16x16_car_red
		449 =>	x"02020202",
		450 =>	x"02020202",
		451 =>	x"02020202",
		452 =>	x"02020000",
		453 =>	x"00020202",
		454 =>	x"02020202",
		455 =>	x"02020202",
		456 =>	x"02020000",
		457 =>	x"00020203",
		458 =>	x"02020202",
		459 =>	x"02020202",
		460 =>	x"02020200",
		461 =>	x"02020203",
		462 =>	x"03020202",
		463 =>	x"02020202",
		464 =>	x"02020303",
		465 =>	x"03030303",
		466 =>	x"03030202",
		467 =>	x"00000002",
		468 =>	x"02000003",
		469 =>	x"03030303",
		470 =>	x"03030303",
		471 =>	x"00000002",
		472 =>	x"02000000",
		473 =>	x"00060606",
		474 =>	x"03030303",
		475 =>	x"02000202",
		476 =>	x"02020303",
		477 =>	x"03060606",
		478 =>	x"06030303",
		479 =>	x"03030302",
		480 =>	x"02020303",
		481 =>	x"03060606",
		482 =>	x"06030303",
		483 =>	x"03030302",
		484 =>	x"02000000",
		485 =>	x"00060606",
		486 =>	x"03030303",
		487 =>	x"02000202",
		488 =>	x"02000003",
		489 =>	x"03030303",
		490 =>	x"03030303",
		491 =>	x"00000002",
		492 =>	x"02020303",
		493 =>	x"03030303",
		494 =>	x"03030202",
		495 =>	x"00000002",
		496 =>	x"02020200",
		497 =>	x"02020203",
		498 =>	x"03020202",
		499 =>	x"02020202",
		500 =>	x"02020000",
		501 =>	x"00020203",
		502 =>	x"02020202",
		503 =>	x"02020202",
		504 =>	x"02020000",
		505 =>	x"00020202",
		506 =>	x"02020202",
		507 =>	x"02020202",
		508 =>	x"02020202",
		509 =>	x"02020202",
		510 =>	x"02020202",
		511 =>	x"02020202",
		512 =>	x"01010101", -- IMG_16x16_flag
		513 =>	x"01010101",
		514 =>	x"01010101",
		515 =>	x"01010101",
		516 =>	x"01010606",
		517 =>	x"01010101",
		518 =>	x"01010101",
		519 =>	x"01010101",
		520 =>	x"01010606",
		521 =>	x"06060101",
		522 =>	x"01010101",
		523 =>	x"01010101",
		524 =>	x"01010606",
		525 =>	x"06060606",
		526 =>	x"01010101",
		527 =>	x"01010101",
		528 =>	x"01010606",
		529 =>	x"06060606",
		530 =>	x"06060101",
		531 =>	x"01010101",
		532 =>	x"01010606",
		533 =>	x"06060606",
		534 =>	x"06060606",
		535 =>	x"01010101",
		536 =>	x"01010606",
		537 =>	x"06060606",
		538 =>	x"06060101",
		539 =>	x"01010101",
		540 =>	x"01010606",
		541 =>	x"06060606",
		542 =>	x"01010101",
		543 =>	x"01010101",
		544 =>	x"01010606",
		545 =>	x"06060101",
		546 =>	x"01010101",
		547 =>	x"01010101",
		548 =>	x"01010606",
		549 =>	x"01010101",
		550 =>	x"01010101",
		551 =>	x"01010101",
		552 =>	x"01010606",
		553 =>	x"01010101",
		554 =>	x"01010101",
		555 =>	x"01010101",
		556 =>	x"01010606",
		557 =>	x"01010101",
		558 =>	x"01010101",
		559 =>	x"01010101",
		560 =>	x"01010606",
		561 =>	x"01010101",
		562 =>	x"01010101",
		563 =>	x"01010101",
		564 =>	x"01060606",
		565 =>	x"06010101",
		566 =>	x"01010101",
		567 =>	x"01010101",
		568 =>	x"01060606",
		569 =>	x"06010101",
		570 =>	x"01010101",
		571 =>	x"01010101",
		572 =>	x"01010101",
		573 =>	x"01010101",
		574 =>	x"01010101",
		575 =>	x"01010101",
		576 =>	x"07070707", -- IMG_16x16_map_element_00
		577 =>	x"07070807",
		578 =>	x"08080707",
		579 =>	x"07070707",
		580 =>	x"07070707",
		581 =>	x"090A0A09",
		582 =>	x"0A090A08",
		583 =>	x"07070707",
		584 =>	x"0707080A",
		585 =>	x"090A0A09",
		586 =>	x"0B0C0A0A",
		587 =>	x"07070707",
		588 =>	x"0707090A",
		589 =>	x"0A0A0909",
		590 =>	x"0A0A0909",
		591 =>	x"0A0A0707",
		592 =>	x"07080A0A",
		593 =>	x"0A0A0909",
		594 =>	x"0A030909",
		595 =>	x"09080807",
		596 =>	x"0809090A",
		597 =>	x"0A030909",
		598 =>	x"0A03090A",
		599 =>	x"0A0A0A08",
		600 =>	x"080A0A0A",
		601 =>	x"0A0A0A09",
		602 =>	x"0A0A0A03",
		603 =>	x"030A0A08",
		604 =>	x"080B0909",
		605 =>	x"0A090908",
		606 =>	x"09090A09",
		607 =>	x"030A0808",
		608 =>	x"080A0A0B",
		609 =>	x"0A0A0A0A",
		610 =>	x"0A0A0A03",
		611 =>	x"0A0A0A08",
		612 =>	x"080A0A0A",
		613 =>	x"0A0B0A09",
		614 =>	x"0A0A090A",
		615 =>	x"090A0908",
		616 =>	x"08090A0A",
		617 =>	x"0A0A090A",
		618 =>	x"03090A0A",
		619 =>	x"09080908",
		620 =>	x"070A0A09",
		621 =>	x"0909090A",
		622 =>	x"0A09090A",
		623 =>	x"09090807",
		624 =>	x"0707090A",
		625 =>	x"0A090A0A",
		626 =>	x"0909090A",
		627 =>	x"0A0A0807",
		628 =>	x"0707080B",
		629 =>	x"0A090B0A",
		630 =>	x"09090A0A",
		631 =>	x"09080707",
		632 =>	x"07070707",
		633 =>	x"080A0B0B",
		634 =>	x"0A030807",
		635 =>	x"07070707",
		636 =>	x"07070707",
		637 =>	x"07070808",
		638 =>	x"08080707",
		639 =>	x"07070707",
		640 =>	x"0D0D0D0D", -- IMG_16x16_map_element_01
		641 =>	x"0D0D0D0D",
		642 =>	x"0D0D0D0D",
		643 =>	x"0D0D0E0F",
		644 =>	x"0D0D0D0D",
		645 =>	x"0D0D0D0D",
		646 =>	x"0D0D0D0D",
		647 =>	x"0D0D0E0F",
		648 =>	x"0D0D0D0D",
		649 =>	x"0D0D0D0D",
		650 =>	x"0D0D0D0D",
		651 =>	x"0D0D0E0F",
		652 =>	x"0D0D0D0D",
		653 =>	x"0D0D0D0D",
		654 =>	x"0D0D0D0D",
		655 =>	x"0D0D0E0F",
		656 =>	x"0D0D0D0D",
		657 =>	x"0D0D0D0D",
		658 =>	x"0D0D0D0D",
		659 =>	x"0D0D0E0F",
		660 =>	x"0D0D0D0D",
		661 =>	x"0D0D0D0D",
		662 =>	x"0D0D0D0D",
		663 =>	x"0D0D0E0F",
		664 =>	x"0D0D0D0D",
		665 =>	x"0D0D0D0D",
		666 =>	x"0D0D0D0D",
		667 =>	x"0D0D0E0F",
		668 =>	x"0D0D0D0D",
		669 =>	x"0D0D0D0D",
		670 =>	x"0D0D0D0D",
		671 =>	x"0D0D0E0F",
		672 =>	x"0D0D0D0D",
		673 =>	x"0D0D0D0D",
		674 =>	x"0D0D0D0D",
		675 =>	x"0D0D0E0F",
		676 =>	x"0D0D0D0D",
		677 =>	x"0D0D0D0D",
		678 =>	x"0D0D0D0D",
		679 =>	x"0D0D0E0F",
		680 =>	x"0D0D0D0D",
		681 =>	x"0D0D0D0D",
		682 =>	x"0D0D0D0D",
		683 =>	x"0D0D0E0F",
		684 =>	x"0D0D0D0D",
		685 =>	x"0D0D0D0D",
		686 =>	x"0D0D0D0D",
		687 =>	x"0D0D0E0F",
		688 =>	x"0D0D0D0D",
		689 =>	x"0D0D0D0D",
		690 =>	x"0D0D0D0D",
		691 =>	x"0D0D0E0F",
		692 =>	x"0D0D0D0D",
		693 =>	x"0D0D0D0D",
		694 =>	x"0D0D0D0D",
		695 =>	x"0D0D0E0F",
		696 =>	x"0D0D0D0D",
		697 =>	x"0D0D0D0D",
		698 =>	x"0D0D0D0D",
		699 =>	x"0D0D0E0F",
		700 =>	x"0D0D0D0D",
		701 =>	x"0D0D0D0D",
		702 =>	x"0D0D0D0D",
		703 =>	x"0D0D0E0F",
		704 =>	x"1011120F", -- IMG_16x16_map_element_02
		705 =>	x"0F0F0F0F",
		706 =>	x"0F0F0F0F",
		707 =>	x"0F0F0F0F",
		708 =>	x"13141516",
		709 =>	x"0E0E0E0E",
		710 =>	x"0E0E0E0E",
		711 =>	x"0E0E0E0E",
		712 =>	x"12170D0D",
		713 =>	x"0D0D0D0D",
		714 =>	x"0D0D0D0D",
		715 =>	x"0D0D0D0D",
		716 =>	x"0F0E0D0D",
		717 =>	x"0D0D0D0D",
		718 =>	x"0D0D0D0D",
		719 =>	x"0D0D0D0D",
		720 =>	x"0F0E0D0D",
		721 =>	x"0D0D0D0D",
		722 =>	x"0D0D0D0D",
		723 =>	x"0D0D0D0D",
		724 =>	x"0F0E0D0D",
		725 =>	x"0D0D0D0D",
		726 =>	x"0D0D0D0D",
		727 =>	x"0D0D0D0D",
		728 =>	x"0F0E0D0D",
		729 =>	x"0D0D0D0D",
		730 =>	x"0D0D0D0D",
		731 =>	x"0D0D0D0D",
		732 =>	x"0F0E0D0D",
		733 =>	x"0D0D0D0D",
		734 =>	x"0D0D0D0D",
		735 =>	x"0D0D0D0D",
		736 =>	x"0F0E0D0D",
		737 =>	x"0D0D0D0D",
		738 =>	x"0D0D0D0D",
		739 =>	x"0D0D0D0D",
		740 =>	x"0F0E0D0D",
		741 =>	x"0D0D0D0D",
		742 =>	x"0D0D0D0D",
		743 =>	x"0D0D0D0D",
		744 =>	x"0F0E0D0D",
		745 =>	x"0D0D0D0D",
		746 =>	x"0D0D0D0D",
		747 =>	x"0D0D0D0D",
		748 =>	x"0F0E0D0D",
		749 =>	x"0D0D0D0D",
		750 =>	x"0D0D0D0D",
		751 =>	x"0D0D0D0D",
		752 =>	x"0F0E0D0D",
		753 =>	x"0D0D0D0D",
		754 =>	x"0D0D0D0D",
		755 =>	x"0D0D0D0D",
		756 =>	x"12170D0D",
		757 =>	x"0D0D0D0D",
		758 =>	x"0D0D0D0D",
		759 =>	x"0D0D0D0D",
		760 =>	x"13141516",
		761 =>	x"0E0E0E0E",
		762 =>	x"0E0E0E0E",
		763 =>	x"0E0E0E0E",
		764 =>	x"1011120F",
		765 =>	x"0F0F0F0F",
		766 =>	x"0F0F0F0F",
		767 =>	x"0F0F0F0F",
		768 =>	x"0F0E0D0D", -- IMG_16x16_map_element_03
		769 =>	x"0D0D0D0D",
		770 =>	x"0D0D0D0D",
		771 =>	x"0D0D0E0F",
		772 =>	x"0E180D0D",
		773 =>	x"0D0D0D0D",
		774 =>	x"0D0D0D0D",
		775 =>	x"0D0D180E",
		776 =>	x"0D0D0D0D",
		777 =>	x"0D0D0D0D",
		778 =>	x"0D0D0D0D",
		779 =>	x"0D0D0D0D",
		780 =>	x"0D0D0D0D",
		781 =>	x"0D0D0D0D",
		782 =>	x"0D0D0D0D",
		783 =>	x"0D0D0D0D",
		784 =>	x"0D0D0D0D",
		785 =>	x"0D0D0D0D",
		786 =>	x"0D0D0D0D",
		787 =>	x"0D0D0D0D",
		788 =>	x"0D0D0D0D",
		789 =>	x"0D0D0D0D",
		790 =>	x"0D0D0D0D",
		791 =>	x"0D0D0D0D",
		792 =>	x"0D0D0D0D",
		793 =>	x"0D0D0D0D",
		794 =>	x"0D0D0D0D",
		795 =>	x"0D0D0D0D",
		796 =>	x"0D0D0D0D",
		797 =>	x"0D0D0D0D",
		798 =>	x"0D0D0D0D",
		799 =>	x"0D0D0D0D",
		800 =>	x"0D0D0D0D",
		801 =>	x"0D0D0D0D",
		802 =>	x"0D0D0D0D",
		803 =>	x"0D0D0D0D",
		804 =>	x"0D0D0D0D",
		805 =>	x"0D0D0D0D",
		806 =>	x"0D0D0D0D",
		807 =>	x"0D0D0D0D",
		808 =>	x"0D0D0D0D",
		809 =>	x"0D0D0D0D",
		810 =>	x"0D0D0D0D",
		811 =>	x"0D0D0D0D",
		812 =>	x"0D0D0D0D",
		813 =>	x"0D0D0D0D",
		814 =>	x"0D0D0D0D",
		815 =>	x"0D0D0D0D",
		816 =>	x"0D0D0D0D",
		817 =>	x"0D0D0D0D",
		818 =>	x"0D0D0D0D",
		819 =>	x"0D0D0D0D",
		820 =>	x"0D0D0D0D",
		821 =>	x"0D0D0D0D",
		822 =>	x"0D0D0D0D",
		823 =>	x"0D0D0D0D",
		824 =>	x"0E180D0D",
		825 =>	x"0D0D0D0D",
		826 =>	x"0D0D0D0D",
		827 =>	x"0D0D180E",
		828 =>	x"0F0E0D0D",
		829 =>	x"0D0D0D0D",
		830 =>	x"0D0D0D0D",
		831 =>	x"0D0D0E0F",
		832 =>	x"0F0F0F0F", -- IMG_16x16_map_element_04
		833 =>	x"0F0F0F0F",
		834 =>	x"0F0F0F0F",
		835 =>	x"0F121110",
		836 =>	x"0E0E0E0E",
		837 =>	x"0E0E0E0E",
		838 =>	x"0E0E0E0E",
		839 =>	x"16151413",
		840 =>	x"0D0D0D0D",
		841 =>	x"0D0D0D0D",
		842 =>	x"0D0D0D0D",
		843 =>	x"0D0D1712",
		844 =>	x"0D0D0D0D",
		845 =>	x"0D0D0D0D",
		846 =>	x"0D0D0D0D",
		847 =>	x"0D0D0E0F",
		848 =>	x"0D0D0D0D",
		849 =>	x"0D0D0D0D",
		850 =>	x"0D0D0D0D",
		851 =>	x"0D0D0E0F",
		852 =>	x"0D0D0D0D",
		853 =>	x"0D0D0D0D",
		854 =>	x"0D0D0D0D",
		855 =>	x"0D0D0E0F",
		856 =>	x"0D0D0D0D",
		857 =>	x"0D0D0D0D",
		858 =>	x"0D0D0D0D",
		859 =>	x"0D0D0E0F",
		860 =>	x"0D0D0D0D",
		861 =>	x"0D0D0D0D",
		862 =>	x"0D0D0D0D",
		863 =>	x"0D0D0E0F",
		864 =>	x"0D0D0D0D",
		865 =>	x"0D0D0D0D",
		866 =>	x"0D0D0D0D",
		867 =>	x"0D0D0E0F",
		868 =>	x"0D0D0D0D",
		869 =>	x"0D0D0D0D",
		870 =>	x"0D0D0D0D",
		871 =>	x"0D0D0E0F",
		872 =>	x"0D0D0D0D",
		873 =>	x"0D0D0D0D",
		874 =>	x"0D0D0D0D",
		875 =>	x"0D0D0E0F",
		876 =>	x"0D0D0D0D",
		877 =>	x"0D0D0D0D",
		878 =>	x"0D0D0D0D",
		879 =>	x"0D0D0E0F",
		880 =>	x"0D0D0D0D",
		881 =>	x"0D0D0D0D",
		882 =>	x"0D0D0D0D",
		883 =>	x"0D0D0E0F",
		884 =>	x"0D0D0D0D",
		885 =>	x"0D0D0D0D",
		886 =>	x"0D0D0D0D",
		887 =>	x"0D0D1712",
		888 =>	x"0E0E0E0E",
		889 =>	x"0E0E0E0E",
		890 =>	x"0E0E0E0E",
		891 =>	x"16151413",
		892 =>	x"0F0F0F0F",
		893 =>	x"0F0F0F0F",
		894 =>	x"0F0F0F0F",
		895 =>	x"0F121110",
		896 =>	x"0F0E0D0D", -- IMG_16x16_map_element_05
		897 =>	x"0D0D0D0D",
		898 =>	x"0D0D0D0D",
		899 =>	x"0D0D0D0D",
		900 =>	x"0F0E0D0D",
		901 =>	x"0D0D0D0D",
		902 =>	x"0D0D0D0D",
		903 =>	x"0D0D0D0D",
		904 =>	x"0F0E0D0D",
		905 =>	x"0D0D0D0D",
		906 =>	x"0D0D0D0D",
		907 =>	x"0D0D0D0D",
		908 =>	x"0F0E0D0D",
		909 =>	x"0D0D0D0D",
		910 =>	x"0D0D0D0D",
		911 =>	x"0D0D0D0D",
		912 =>	x"0F0E0D0D",
		913 =>	x"0D0D0D0D",
		914 =>	x"0D0D0D0D",
		915 =>	x"0D0D0D0D",
		916 =>	x"0F0E0D0D",
		917 =>	x"0D0D0D0D",
		918 =>	x"0D0D0D0D",
		919 =>	x"0D0D0D0D",
		920 =>	x"0F0E0D0D",
		921 =>	x"0D0D0D0D",
		922 =>	x"0D0D0D0D",
		923 =>	x"0D0D0D0D",
		924 =>	x"0F0E0D0D",
		925 =>	x"0D0D0D0D",
		926 =>	x"0D0D0D0D",
		927 =>	x"0D0D0D0D",
		928 =>	x"0F0E0D0D",
		929 =>	x"0D0D0D0D",
		930 =>	x"0D0D0D0D",
		931 =>	x"0D0D0D0D",
		932 =>	x"0F0E0D0D",
		933 =>	x"0D0D0D0D",
		934 =>	x"0D0D0D0D",
		935 =>	x"0D0D0D0D",
		936 =>	x"0F0E0D0D",
		937 =>	x"0D0D0D0D",
		938 =>	x"0D0D0D0D",
		939 =>	x"0D0D0D0D",
		940 =>	x"0F0E0D0D",
		941 =>	x"0D0D0D0D",
		942 =>	x"0D0D0D0D",
		943 =>	x"0D0D0D0D",
		944 =>	x"0F0E0D0D",
		945 =>	x"0D0D0D0D",
		946 =>	x"0D0D0D0D",
		947 =>	x"0D0D0D0D",
		948 =>	x"12170D0D",
		949 =>	x"0D0D0D0D",
		950 =>	x"0D0D0D0D",
		951 =>	x"0D0D0D0D",
		952 =>	x"13141516",
		953 =>	x"0E0E0E0E",
		954 =>	x"0E0E0E0E",
		955 =>	x"0E0E0E0E",
		956 =>	x"1011120F",
		957 =>	x"0F0F0F0F",
		958 =>	x"0F0F0F0F",
		959 =>	x"0F0F0F0F",
		960 =>	x"0D0D0D0D", -- IMG_16x16_map_element_06
		961 =>	x"0D0D0D0D",
		962 =>	x"0D0D0D0D",
		963 =>	x"0D0D0D0D",
		964 =>	x"0D0D0D0D",
		965 =>	x"0D0D0D0D",
		966 =>	x"0D0D0D0D",
		967 =>	x"0D0D0D0D",
		968 =>	x"0D0D0D0D",
		969 =>	x"0D0D0D0D",
		970 =>	x"0D0D0D0D",
		971 =>	x"0D0D0D0D",
		972 =>	x"0D0D0D0D",
		973 =>	x"0D0D0D0D",
		974 =>	x"0D0D0D0D",
		975 =>	x"0D0D0D0D",
		976 =>	x"0D0D0D0D",
		977 =>	x"0D0D0D0D",
		978 =>	x"0D0D0D0D",
		979 =>	x"0D0D0D0D",
		980 =>	x"0D0D0D0D",
		981 =>	x"0D0D0D0D",
		982 =>	x"0D0D0D0D",
		983 =>	x"0D0D0D0D",
		984 =>	x"0D0D0D0D",
		985 =>	x"0D0D0D0D",
		986 =>	x"0D0D0D0D",
		987 =>	x"0D0D0D0D",
		988 =>	x"0D0D0D0D",
		989 =>	x"0D0D0D0D",
		990 =>	x"0D0D0D0D",
		991 =>	x"0D0D0D0D",
		992 =>	x"0D0D0D0D",
		993 =>	x"0D0D0D0D",
		994 =>	x"0D0D0D0D",
		995 =>	x"0D0D0D0D",
		996 =>	x"0D0D0D0D",
		997 =>	x"0D0D0D0D",
		998 =>	x"0D0D0D0D",
		999 =>	x"0D0D0D0D",
		1000 =>	x"0D0D0D0D",
		1001 =>	x"0D0D0D0D",
		1002 =>	x"0D0D0D0D",
		1003 =>	x"0D0D0D0D",
		1004 =>	x"0D0D0D0D",
		1005 =>	x"0D0D0D0D",
		1006 =>	x"0D0D0D0D",
		1007 =>	x"0D0D0D0D",
		1008 =>	x"0D0D0D0D",
		1009 =>	x"0D0D0D0D",
		1010 =>	x"0D0D0D0D",
		1011 =>	x"0D0D0D0D",
		1012 =>	x"0D0D0D0D",
		1013 =>	x"0D0D0D0D",
		1014 =>	x"0D0D0D0D",
		1015 =>	x"0D0D0D0D",
		1016 =>	x"0E0E0E0E",
		1017 =>	x"0E0E0E0E",
		1018 =>	x"0E0E0E0E",
		1019 =>	x"0E0E0E0E",
		1020 =>	x"0F0F0F0F",
		1021 =>	x"0F0F0F0F",
		1022 =>	x"0F0F0F0F",
		1023 =>	x"0F0F0F0F",
		1024 =>	x"0D0D0D0D", -- IMG_16x16_map_element_07
		1025 =>	x"0D0D0D0D",
		1026 =>	x"0D0D0D0D",
		1027 =>	x"0D0D0E0F",
		1028 =>	x"0D0D0D0D",
		1029 =>	x"0D0D0D0D",
		1030 =>	x"0D0D0D0D",
		1031 =>	x"0D0D0E0F",
		1032 =>	x"0D0D0D0D",
		1033 =>	x"0D0D0D0D",
		1034 =>	x"0D0D0D0D",
		1035 =>	x"0D0D0E0F",
		1036 =>	x"0D0D0D0D",
		1037 =>	x"0D0D0D0D",
		1038 =>	x"0D0D0D0D",
		1039 =>	x"0D0D0E0F",
		1040 =>	x"0D0D0D0D",
		1041 =>	x"0D0D0D0D",
		1042 =>	x"0D0D0D0D",
		1043 =>	x"0D0D0E0F",
		1044 =>	x"0D0D0D0D",
		1045 =>	x"0D0D0D0D",
		1046 =>	x"0D0D0D0D",
		1047 =>	x"0D0D0E0F",
		1048 =>	x"0D0D0D0D",
		1049 =>	x"0D0D0D0D",
		1050 =>	x"0D0D0D0D",
		1051 =>	x"0D0D0E0F",
		1052 =>	x"0D0D0D0D",
		1053 =>	x"0D0D0D0D",
		1054 =>	x"0D0D0D0D",
		1055 =>	x"0D0D0E0F",
		1056 =>	x"0D0D0D0D",
		1057 =>	x"0D0D0D0D",
		1058 =>	x"0D0D0D0D",
		1059 =>	x"0D0D0E0F",
		1060 =>	x"0D0D0D0D",
		1061 =>	x"0D0D0D0D",
		1062 =>	x"0D0D0D0D",
		1063 =>	x"0D0D0E0F",
		1064 =>	x"0D0D0D0D",
		1065 =>	x"0D0D0D0D",
		1066 =>	x"0D0D0D0D",
		1067 =>	x"0D0D0E0F",
		1068 =>	x"0D0D0D0D",
		1069 =>	x"0D0D0D0D",
		1070 =>	x"0D0D0D0D",
		1071 =>	x"0D0D0E0F",
		1072 =>	x"0D0D0D0D",
		1073 =>	x"0D0D0D0D",
		1074 =>	x"0D0D0D0D",
		1075 =>	x"0D0D0E0F",
		1076 =>	x"0D0D0D0D",
		1077 =>	x"0D0D0D0D",
		1078 =>	x"0D0D0D0D",
		1079 =>	x"0D0D1712",
		1080 =>	x"0E0E0E0E",
		1081 =>	x"0E0E0E0E",
		1082 =>	x"0E0E0E0E",
		1083 =>	x"16151413",
		1084 =>	x"0F0F0F0F",
		1085 =>	x"0F0F0F0F",
		1086 =>	x"0F0F0F0F",
		1087 =>	x"0F121110",
		1088 =>	x"0F0E0D0D", -- IMG_16x16_map_element_08
		1089 =>	x"0D0D0D0D",
		1090 =>	x"0D0D0D0D",
		1091 =>	x"0D0D0E0F",
		1092 =>	x"0F0E0D0D",
		1093 =>	x"0D0D0D0D",
		1094 =>	x"0D0D0D0D",
		1095 =>	x"0D0D180E",
		1096 =>	x"0F0E0D0D",
		1097 =>	x"0D0D0D0D",
		1098 =>	x"0D0D0D0D",
		1099 =>	x"0D0D0D0D",
		1100 =>	x"0F0E0D0D",
		1101 =>	x"0D0D0D0D",
		1102 =>	x"0D0D0D0D",
		1103 =>	x"0D0D0D0D",
		1104 =>	x"0F0E0D0D",
		1105 =>	x"0D0D0D0D",
		1106 =>	x"0D0D0D0D",
		1107 =>	x"0D0D0D0D",
		1108 =>	x"0F0E0D0D",
		1109 =>	x"0D0D0D0D",
		1110 =>	x"0D0D0D0D",
		1111 =>	x"0D0D0D0D",
		1112 =>	x"0F0E0D0D",
		1113 =>	x"0D0D0D0D",
		1114 =>	x"0D0D0D0D",
		1115 =>	x"0D0D0D0D",
		1116 =>	x"0F0E0D0D",
		1117 =>	x"0D0D0D0D",
		1118 =>	x"0D0D0D0D",
		1119 =>	x"0D0D0D0D",
		1120 =>	x"0F0E0D0D",
		1121 =>	x"0D0D0D0D",
		1122 =>	x"0D0D0D0D",
		1123 =>	x"0D0D0D0D",
		1124 =>	x"0F0E0D0D",
		1125 =>	x"0D0D0D0D",
		1126 =>	x"0D0D0D0D",
		1127 =>	x"0D0D0D0D",
		1128 =>	x"0F0E0D0D",
		1129 =>	x"0D0D0D0D",
		1130 =>	x"0D0D0D0D",
		1131 =>	x"0D0D0D0D",
		1132 =>	x"0F0E0D0D",
		1133 =>	x"0D0D0D0D",
		1134 =>	x"0D0D0D0D",
		1135 =>	x"0D0D0D0D",
		1136 =>	x"0F0E0D0D",
		1137 =>	x"0D0D0D0D",
		1138 =>	x"0D0D0D0D",
		1139 =>	x"0D0D0D0D",
		1140 =>	x"12170D0D",
		1141 =>	x"0D0D0D0D",
		1142 =>	x"0D0D0D0D",
		1143 =>	x"0D0D0D0D",
		1144 =>	x"13141516",
		1145 =>	x"0E0E0E0E",
		1146 =>	x"0E0E0E0E",
		1147 =>	x"0E0E0E0E",
		1148 =>	x"1011120F",
		1149 =>	x"0F0F0F0F",
		1150 =>	x"0F0F0F0F",
		1151 =>	x"0F0F0F0F",
		1152 =>	x"0F0E0D0D", -- IMG_16x16_map_element_09
		1153 =>	x"0D0D0D0D",
		1154 =>	x"0D0D0D0D",
		1155 =>	x"0D0D0E0F",
		1156 =>	x"0F0E0D0D",
		1157 =>	x"0D0D0D0D",
		1158 =>	x"0D0D0D0D",
		1159 =>	x"0D0D0E0F",
		1160 =>	x"0F0E0D0D",
		1161 =>	x"0D0D0D0D",
		1162 =>	x"0D0D0D0D",
		1163 =>	x"0D0D0E0F",
		1164 =>	x"0F0E0D0D",
		1165 =>	x"0D0D0D0D",
		1166 =>	x"0D0D0D0D",
		1167 =>	x"0D0D0E0F",
		1168 =>	x"0F0E0D0D",
		1169 =>	x"0D0D0D0D",
		1170 =>	x"0D0D0D0D",
		1171 =>	x"0D0D0E0F",
		1172 =>	x"0F0E0D0D",
		1173 =>	x"0D0D0D0D",
		1174 =>	x"0D0D0D0D",
		1175 =>	x"0D0D0E0F",
		1176 =>	x"0F0E0D0D",
		1177 =>	x"0D0D0D0D",
		1178 =>	x"0D0D0D0D",
		1179 =>	x"0D0D0E0F",
		1180 =>	x"0F0E0D0D",
		1181 =>	x"0D0D0D0D",
		1182 =>	x"0D0D0D0D",
		1183 =>	x"0D0D0E0F",
		1184 =>	x"0F0E0D0D",
		1185 =>	x"0D0D0D0D",
		1186 =>	x"0D0D0D0D",
		1187 =>	x"0D0D0E0F",
		1188 =>	x"0F0E0D0D",
		1189 =>	x"0D0D0D0D",
		1190 =>	x"0D0D0D0D",
		1191 =>	x"0D0D0E0F",
		1192 =>	x"0F0E0D0D",
		1193 =>	x"0D0D0D0D",
		1194 =>	x"0D0D0D0D",
		1195 =>	x"0D0D0E0F",
		1196 =>	x"0F0E0D0D",
		1197 =>	x"0D0D0D0D",
		1198 =>	x"0D0D0D0D",
		1199 =>	x"0D0D0E0F",
		1200 =>	x"0F0E0D0D",
		1201 =>	x"0D0D0D0D",
		1202 =>	x"0D0D0D0D",
		1203 =>	x"0D0D0E0F",
		1204 =>	x"12170D0D",
		1205 =>	x"0D0D0D0D",
		1206 =>	x"0D0D0D0D",
		1207 =>	x"0D0D1712",
		1208 =>	x"13141516",
		1209 =>	x"0E0E0E0E",
		1210 =>	x"0E0E0E0E",
		1211 =>	x"16151413",
		1212 =>	x"1011120F",
		1213 =>	x"0F0F0F0F",
		1214 =>	x"0F0F0F0F",
		1215 =>	x"0F121110",
		1216 =>	x"0F0E0D0D", -- IMG_16x16_map_element_10
		1217 =>	x"0D0D0D0D",
		1218 =>	x"0D0D0D0D",
		1219 =>	x"0D0D0E0F",
		1220 =>	x"0E180D0D",
		1221 =>	x"0D0D0D0D",
		1222 =>	x"0D0D0D0D",
		1223 =>	x"0D0D0E0F",
		1224 =>	x"0D0D0D0D",
		1225 =>	x"0D0D0D0D",
		1226 =>	x"0D0D0D0D",
		1227 =>	x"0D0D0E0F",
		1228 =>	x"0D0D0D0D",
		1229 =>	x"0D0D0D0D",
		1230 =>	x"0D0D0D0D",
		1231 =>	x"0D0D0E0F",
		1232 =>	x"0D0D0D0D",
		1233 =>	x"0D0D0D0D",
		1234 =>	x"0D0D0D0D",
		1235 =>	x"0D0D0E0F",
		1236 =>	x"0D0D0D0D",
		1237 =>	x"0D0D0D0D",
		1238 =>	x"0D0D0D0D",
		1239 =>	x"0D0D0E0F",
		1240 =>	x"0D0D0D0D",
		1241 =>	x"0D0D0D0D",
		1242 =>	x"0D0D0D0D",
		1243 =>	x"0D0D0E0F",
		1244 =>	x"0D0D0D0D",
		1245 =>	x"0D0D0D0D",
		1246 =>	x"0D0D0D0D",
		1247 =>	x"0D0D0E0F",
		1248 =>	x"0D0D0D0D",
		1249 =>	x"0D0D0D0D",
		1250 =>	x"0D0D0D0D",
		1251 =>	x"0D0D0E0F",
		1252 =>	x"0D0D0D0D",
		1253 =>	x"0D0D0D0D",
		1254 =>	x"0D0D0D0D",
		1255 =>	x"0D0D0E0F",
		1256 =>	x"0D0D0D0D",
		1257 =>	x"0D0D0D0D",
		1258 =>	x"0D0D0D0D",
		1259 =>	x"0D0D0E0F",
		1260 =>	x"0D0D0D0D",
		1261 =>	x"0D0D0D0D",
		1262 =>	x"0D0D0D0D",
		1263 =>	x"0D0D0E0F",
		1264 =>	x"0D0D0D0D",
		1265 =>	x"0D0D0D0D",
		1266 =>	x"0D0D0D0D",
		1267 =>	x"0D0D0E0F",
		1268 =>	x"0D0D0D0D",
		1269 =>	x"0D0D0D0D",
		1270 =>	x"0D0D0D0D",
		1271 =>	x"0D0D1712",
		1272 =>	x"0E0E0E0E",
		1273 =>	x"0E0E0E0E",
		1274 =>	x"0E0E0E0E",
		1275 =>	x"16151413",
		1276 =>	x"0F0F0F0F",
		1277 =>	x"0F0F0F0F",
		1278 =>	x"0F0F0F0F",
		1279 =>	x"0F121110",
		1280 =>	x"1011120F", -- IMG_16x16_map_element_11
		1281 =>	x"0F0F0F0F",
		1282 =>	x"0F0F0F0F",
		1283 =>	x"0F0F0F0F",
		1284 =>	x"13141516",
		1285 =>	x"0E0E0E0E",
		1286 =>	x"0E0E0E0E",
		1287 =>	x"0E0E0E0E",
		1288 =>	x"12170D0D",
		1289 =>	x"0D0D0D0D",
		1290 =>	x"0D0D0D0D",
		1291 =>	x"0D0D0D0D",
		1292 =>	x"0F0E0D0D",
		1293 =>	x"0D0D0D0D",
		1294 =>	x"0D0D0D0D",
		1295 =>	x"0D0D0D0D",
		1296 =>	x"0F0E0D0D",
		1297 =>	x"0D0D0D0D",
		1298 =>	x"0D0D0D0D",
		1299 =>	x"0D0D0D0D",
		1300 =>	x"0F0E0D0D",
		1301 =>	x"0D0D0D0D",
		1302 =>	x"0D0D0D0D",
		1303 =>	x"0D0D0D0D",
		1304 =>	x"0F0E0D0D",
		1305 =>	x"0D0D0D0D",
		1306 =>	x"0D0D0D0D",
		1307 =>	x"0D0D0D0D",
		1308 =>	x"0F0E0D0D",
		1309 =>	x"0D0D0D0D",
		1310 =>	x"0D0D0D0D",
		1311 =>	x"0D0D0D0D",
		1312 =>	x"0F0E0D0D",
		1313 =>	x"0D0D0D0D",
		1314 =>	x"0D0D0D0D",
		1315 =>	x"0D0D0D0D",
		1316 =>	x"0F0E0D0D",
		1317 =>	x"0D0D0D0D",
		1318 =>	x"0D0D0D0D",
		1319 =>	x"0D0D0D0D",
		1320 =>	x"0F0E0D0D",
		1321 =>	x"0D0D0D0D",
		1322 =>	x"0D0D0D0D",
		1323 =>	x"0D0D0D0D",
		1324 =>	x"0F0E0D0D",
		1325 =>	x"0D0D0D0D",
		1326 =>	x"0D0D0D0D",
		1327 =>	x"0D0D0D0D",
		1328 =>	x"0F0E0D0D",
		1329 =>	x"0D0D0D0D",
		1330 =>	x"0D0D0D0D",
		1331 =>	x"0D0D0D0D",
		1332 =>	x"0F0E0D0D",
		1333 =>	x"0D0D0D0D",
		1334 =>	x"0D0D0D0D",
		1335 =>	x"0D0D0D0D",
		1336 =>	x"0F0E0D0D",
		1337 =>	x"0D0D0D0D",
		1338 =>	x"0D0D0D0D",
		1339 =>	x"0D0D0D0D",
		1340 =>	x"0F0E0D0D",
		1341 =>	x"0D0D0D0D",
		1342 =>	x"0D0D0D0D",
		1343 =>	x"0D0D0D0D",
		1344 =>	x"0F0F0F0F", -- IMG_16x16_map_element_12
		1345 =>	x"0F0F0F0F",
		1346 =>	x"0F0F0F0F",
		1347 =>	x"0F0F0F0F",
		1348 =>	x"0E0E0E0E",
		1349 =>	x"0E0E0E0E",
		1350 =>	x"0E0E0E0E",
		1351 =>	x"0E0E0E0E",
		1352 =>	x"0D0D0D0D",
		1353 =>	x"0D0D0D0D",
		1354 =>	x"0D0D0D0D",
		1355 =>	x"0D0D0D0D",
		1356 =>	x"0D0D0D0D",
		1357 =>	x"0D0D0D0D",
		1358 =>	x"0D0D0D0D",
		1359 =>	x"0D0D0D0D",
		1360 =>	x"0D0D0D0D",
		1361 =>	x"0D0D0D0D",
		1362 =>	x"0D0D0D0D",
		1363 =>	x"0D0D0D0D",
		1364 =>	x"0D0D0D0D",
		1365 =>	x"0D0D0D0D",
		1366 =>	x"0D0D0D0D",
		1367 =>	x"0D0D0D0D",
		1368 =>	x"0D0D0D0D",
		1369 =>	x"0D0D0D0D",
		1370 =>	x"0D0D0D0D",
		1371 =>	x"0D0D0D0D",
		1372 =>	x"0D0D0D0D",
		1373 =>	x"0D0D0D0D",
		1374 =>	x"0D0D0D0D",
		1375 =>	x"0D0D0D0D",
		1376 =>	x"0D0D0D0D",
		1377 =>	x"0D0D0D0D",
		1378 =>	x"0D0D0D0D",
		1379 =>	x"0D0D0D0D",
		1380 =>	x"0D0D0D0D",
		1381 =>	x"0D0D0D0D",
		1382 =>	x"0D0D0D0D",
		1383 =>	x"0D0D0D0D",
		1384 =>	x"0D0D0D0D",
		1385 =>	x"0D0D0D0D",
		1386 =>	x"0D0D0D0D",
		1387 =>	x"0D0D0D0D",
		1388 =>	x"0D0D0D0D",
		1389 =>	x"0D0D0D0D",
		1390 =>	x"0D0D0D0D",
		1391 =>	x"0D0D0D0D",
		1392 =>	x"0D0D0D0D",
		1393 =>	x"0D0D0D0D",
		1394 =>	x"0D0D0D0D",
		1395 =>	x"0D0D0D0D",
		1396 =>	x"0D0D0D0D",
		1397 =>	x"0D0D0D0D",
		1398 =>	x"0D0D0D0D",
		1399 =>	x"0D0D0D0D",
		1400 =>	x"0E180D0D",
		1401 =>	x"0D0D0D0D",
		1402 =>	x"0D0D0D0D",
		1403 =>	x"0D0D180E",
		1404 =>	x"0F0E0D0D",
		1405 =>	x"0D0D0D0D",
		1406 =>	x"0D0D0D0D",
		1407 =>	x"0D0D0E0F",
		1408 =>	x"0F0E0D0D", -- IMG_16x16_map_element_13
		1409 =>	x"0D0D0D0D",
		1410 =>	x"0D0D0D0D",
		1411 =>	x"0D0D0E0F",
		1412 =>	x"0F0E0D0D",
		1413 =>	x"0D0D0D0D",
		1414 =>	x"0D0D0D0D",
		1415 =>	x"0D0D180E",
		1416 =>	x"0F0E0D0D",
		1417 =>	x"0D0D0D0D",
		1418 =>	x"0D0D0D0D",
		1419 =>	x"0D0D0D0D",
		1420 =>	x"0F0E0D0D",
		1421 =>	x"0D0D0D0D",
		1422 =>	x"0D0D0D0D",
		1423 =>	x"0D0D0D0D",
		1424 =>	x"0F0E0D0D",
		1425 =>	x"0D0D0D0D",
		1426 =>	x"0D0D0D0D",
		1427 =>	x"0D0D0D0D",
		1428 =>	x"0F0E0D0D",
		1429 =>	x"0D0D0D0D",
		1430 =>	x"0D0D0D0D",
		1431 =>	x"0D0D0D0D",
		1432 =>	x"0F0E0D0D",
		1433 =>	x"0D0D0D0D",
		1434 =>	x"0D0D0D0D",
		1435 =>	x"0D0D0D0D",
		1436 =>	x"0F0E0D0D",
		1437 =>	x"0D0D0D0D",
		1438 =>	x"0D0D0D0D",
		1439 =>	x"0D0D0D0D",
		1440 =>	x"0F0E0D0D",
		1441 =>	x"0D0D0D0D",
		1442 =>	x"0D0D0D0D",
		1443 =>	x"0D0D0D0D",
		1444 =>	x"0F0E0D0D",
		1445 =>	x"0D0D0D0D",
		1446 =>	x"0D0D0D0D",
		1447 =>	x"0D0D0D0D",
		1448 =>	x"0F0E0D0D",
		1449 =>	x"0D0D0D0D",
		1450 =>	x"0D0D0D0D",
		1451 =>	x"0D0D0D0D",
		1452 =>	x"0F0E0D0D",
		1453 =>	x"0D0D0D0D",
		1454 =>	x"0D0D0D0D",
		1455 =>	x"0D0D0D0D",
		1456 =>	x"0F0E0D0D",
		1457 =>	x"0D0D0D0D",
		1458 =>	x"0D0D0D0D",
		1459 =>	x"0D0D0D0D",
		1460 =>	x"0F0E0D0D",
		1461 =>	x"0D0D0D0D",
		1462 =>	x"0D0D0D0D",
		1463 =>	x"0D0D0D0D",
		1464 =>	x"0F0E0D0D",
		1465 =>	x"0D0D0D0D",
		1466 =>	x"0D0D0D0D",
		1467 =>	x"0D0D180E",
		1468 =>	x"0F0E0D0D",
		1469 =>	x"0D0D0D0D",
		1470 =>	x"0D0D0D0D",
		1471 =>	x"0D0D0E0F",
		1472 =>	x"0F0E0D0D", -- IMG_16x16_map_element_14
		1473 =>	x"0D0D0D0D",
		1474 =>	x"0D0D0D0D",
		1475 =>	x"0D0D0E0F",
		1476 =>	x"0E180D0D",
		1477 =>	x"0D0D0D0D",
		1478 =>	x"0D0D0D0D",
		1479 =>	x"0D0D180E",
		1480 =>	x"0D0D0D0D",
		1481 =>	x"0D0D0D0D",
		1482 =>	x"0D0D0D0D",
		1483 =>	x"0D0D0D0D",
		1484 =>	x"0D0D0D0D",
		1485 =>	x"0D0D0D0D",
		1486 =>	x"0D0D0D0D",
		1487 =>	x"0D0D0D0D",
		1488 =>	x"0D0D0D0D",
		1489 =>	x"0D0D0D0D",
		1490 =>	x"0D0D0D0D",
		1491 =>	x"0D0D0D0D",
		1492 =>	x"0D0D0D0D",
		1493 =>	x"0D0D0D0D",
		1494 =>	x"0D0D0D0D",
		1495 =>	x"0D0D0D0D",
		1496 =>	x"0D0D0D0D",
		1497 =>	x"0D0D0D0D",
		1498 =>	x"0D0D0D0D",
		1499 =>	x"0D0D0D0D",
		1500 =>	x"0D0D0D0D",
		1501 =>	x"0D0D0D0D",
		1502 =>	x"0D0D0D0D",
		1503 =>	x"0D0D0D0D",
		1504 =>	x"0D0D0D0D",
		1505 =>	x"0D0D0D0D",
		1506 =>	x"0D0D0D0D",
		1507 =>	x"0D0D0D0D",
		1508 =>	x"0D0D0D0D",
		1509 =>	x"0D0D0D0D",
		1510 =>	x"0D0D0D0D",
		1511 =>	x"0D0D0D0D",
		1512 =>	x"0D0D0D0D",
		1513 =>	x"0D0D0D0D",
		1514 =>	x"0D0D0D0D",
		1515 =>	x"0D0D0D0D",
		1516 =>	x"0D0D0D0D",
		1517 =>	x"0D0D0D0D",
		1518 =>	x"0D0D0D0D",
		1519 =>	x"0D0D0D0D",
		1520 =>	x"0D0D0D0D",
		1521 =>	x"0D0D0D0D",
		1522 =>	x"0D0D0D0D",
		1523 =>	x"0D0D0D0D",
		1524 =>	x"0D0D0D0D",
		1525 =>	x"0D0D0D0D",
		1526 =>	x"0D0D0D0D",
		1527 =>	x"0D0D0D0D",
		1528 =>	x"0E0E0E0E",
		1529 =>	x"0E0E0E0E",
		1530 =>	x"0E0E0E0E",
		1531 =>	x"0E0E0E0E",
		1532 =>	x"0F0F0F0F",
		1533 =>	x"0F0F0F0F",
		1534 =>	x"0F0F0F0F",
		1535 =>	x"0F0F0F0F",
		1536 =>	x"0F0E0D0D", -- IMG_16x16_map_element_15
		1537 =>	x"0D0D0D0D",
		1538 =>	x"0D0D0D0D",
		1539 =>	x"0D0D0E0F",
		1540 =>	x"0E180D0D",
		1541 =>	x"0D0D0D0D",
		1542 =>	x"0D0D0D0D",
		1543 =>	x"0D0D0E0F",
		1544 =>	x"0D0D0D0D",
		1545 =>	x"0D0D0D0D",
		1546 =>	x"0D0D0D0D",
		1547 =>	x"0D0D0E0F",
		1548 =>	x"0D0D0D0D",
		1549 =>	x"0D0D0D0D",
		1550 =>	x"0D0D0D0D",
		1551 =>	x"0D0D0E0F",
		1552 =>	x"0D0D0D0D",
		1553 =>	x"0D0D0D0D",
		1554 =>	x"0D0D0D0D",
		1555 =>	x"0D0D0E0F",
		1556 =>	x"0D0D0D0D",
		1557 =>	x"0D0D0D0D",
		1558 =>	x"0D0D0D0D",
		1559 =>	x"0D0D0E0F",
		1560 =>	x"0D0D0D0D",
		1561 =>	x"0D0D0D0D",
		1562 =>	x"0D0D0D0D",
		1563 =>	x"0D0D0E0F",
		1564 =>	x"0D0D0D0D",
		1565 =>	x"0D0D0D0D",
		1566 =>	x"0D0D0D0D",
		1567 =>	x"0D0D0E0F",
		1568 =>	x"0D0D0D0D",
		1569 =>	x"0D0D0D0D",
		1570 =>	x"0D0D0D0D",
		1571 =>	x"0D0D0E0F",
		1572 =>	x"0D0D0D0D",
		1573 =>	x"0D0D0D0D",
		1574 =>	x"0D0D0D0D",
		1575 =>	x"0D0D0E0F",
		1576 =>	x"0D0D0D0D",
		1577 =>	x"0D0D0D0D",
		1578 =>	x"0D0D0D0D",
		1579 =>	x"0D0D0E0F",
		1580 =>	x"0D0D0D0D",
		1581 =>	x"0D0D0D0D",
		1582 =>	x"0D0D0D0D",
		1583 =>	x"0D0D0E0F",
		1584 =>	x"0D0D0D0D",
		1585 =>	x"0D0D0D0D",
		1586 =>	x"0D0D0D0D",
		1587 =>	x"0D0D0E0F",
		1588 =>	x"0D0D0D0D",
		1589 =>	x"0D0D0D0D",
		1590 =>	x"0D0D0D0D",
		1591 =>	x"0D0D0E0F",
		1592 =>	x"0E180D0D",
		1593 =>	x"0D0D0D0D",
		1594 =>	x"0D0D0D0D",
		1595 =>	x"0D0D0E0F",
		1596 =>	x"0F0E0D0D",
		1597 =>	x"0D0D0D0D",
		1598 =>	x"0D0D0D0D",
		1599 =>	x"0D0D0E0F",
		1600 =>	x"0F0E0D0D", -- IMG_16x16_map_element_16
		1601 =>	x"0D0D0D0D",
		1602 =>	x"0D0D0D0D",
		1603 =>	x"0D0D0E0F",
		1604 =>	x"0F0E0D0D",
		1605 =>	x"0D0D0D0D",
		1606 =>	x"0D0D0D0D",
		1607 =>	x"0D0D0E0F",
		1608 =>	x"0F0E0D0D",
		1609 =>	x"0D0D0D0D",
		1610 =>	x"0D0D0D0D",
		1611 =>	x"0D0D0E0F",
		1612 =>	x"0F0E0D0D",
		1613 =>	x"0D0D0D0D",
		1614 =>	x"0D0D0D0D",
		1615 =>	x"0D0D0E0F",
		1616 =>	x"0F0E0D0D",
		1617 =>	x"0D0D0D0D",
		1618 =>	x"0D0D0D0D",
		1619 =>	x"0D0D0E0F",
		1620 =>	x"0F0E0D0D",
		1621 =>	x"0D0D0D0D",
		1622 =>	x"0D0D0D0D",
		1623 =>	x"0D0D0E0F",
		1624 =>	x"0F0E0D0D",
		1625 =>	x"0D0D0D0D",
		1626 =>	x"0D0D0D0D",
		1627 =>	x"0D0D0E0F",
		1628 =>	x"0F0E0D0D",
		1629 =>	x"0D0D0D0D",
		1630 =>	x"0D0D0D0D",
		1631 =>	x"0D0D0E0F",
		1632 =>	x"0F0E0D0D",
		1633 =>	x"0D0D0D0D",
		1634 =>	x"0D0D0D0D",
		1635 =>	x"0D0D0E0F",
		1636 =>	x"0F0E0D0D",
		1637 =>	x"0D0D0D0D",
		1638 =>	x"0D0D0D0D",
		1639 =>	x"0D0D0E0F",
		1640 =>	x"0F0E0D0D",
		1641 =>	x"0D0D0D0D",
		1642 =>	x"0D0D0D0D",
		1643 =>	x"0D0D0E0F",
		1644 =>	x"0F0E0D0D",
		1645 =>	x"0D0D0D0D",
		1646 =>	x"0D0D0D0D",
		1647 =>	x"0D0D0E0F",
		1648 =>	x"0F0E0D0D",
		1649 =>	x"0D0D0D0D",
		1650 =>	x"0D0D0D0D",
		1651 =>	x"0D0D0E0F",
		1652 =>	x"0F0E0D0D",
		1653 =>	x"0D0D0D0D",
		1654 =>	x"0D0D0D0D",
		1655 =>	x"0D0D0E0F",
		1656 =>	x"0F0E0D0D",
		1657 =>	x"0D0D0D0D",
		1658 =>	x"0D0D0D0D",
		1659 =>	x"0D0D0E0F",
		1660 =>	x"0F0E0D0D",
		1661 =>	x"0D0D0D0D",
		1662 =>	x"0D0D0D0D",
		1663 =>	x"0D0D0E0F",
		1664 =>	x"0F0F0F0F", -- IMG_16x16_map_element_17
		1665 =>	x"0F0F0F0F",
		1666 =>	x"0F0F0F0F",
		1667 =>	x"0F0F0F0F",
		1668 =>	x"0E0E0E0E",
		1669 =>	x"0E0E0E0E",
		1670 =>	x"0E0E0E0E",
		1671 =>	x"0E0E0E0E",
		1672 =>	x"0D0D0D0D",
		1673 =>	x"0D0D0D0D",
		1674 =>	x"0D0D0D0D",
		1675 =>	x"0D0D0D0D",
		1676 =>	x"0D0D0D0D",
		1677 =>	x"0D0D0D0D",
		1678 =>	x"0D0D0D0D",
		1679 =>	x"0D0D0D0D",
		1680 =>	x"0D0D0D0D",
		1681 =>	x"0D0D0D0D",
		1682 =>	x"0D0D0D0D",
		1683 =>	x"0D0D0D0D",
		1684 =>	x"0D0D0D0D",
		1685 =>	x"0D0D0D0D",
		1686 =>	x"0D0D0D0D",
		1687 =>	x"0D0D0D0D",
		1688 =>	x"0D0D0D0D",
		1689 =>	x"0D0D0D0D",
		1690 =>	x"0D0D0D0D",
		1691 =>	x"0D0D0D0D",
		1692 =>	x"0D0D0D0D",
		1693 =>	x"0D0D0D0D",
		1694 =>	x"0D0D0D0D",
		1695 =>	x"0D0D0D0D",
		1696 =>	x"0D0D0D0D",
		1697 =>	x"0D0D0D0D",
		1698 =>	x"0D0D0D0D",
		1699 =>	x"0D0D0D0D",
		1700 =>	x"0D0D0D0D",
		1701 =>	x"0D0D0D0D",
		1702 =>	x"0D0D0D0D",
		1703 =>	x"0D0D0D0D",
		1704 =>	x"0D0D0D0D",
		1705 =>	x"0D0D0D0D",
		1706 =>	x"0D0D0D0D",
		1707 =>	x"0D0D0D0D",
		1708 =>	x"0D0D0D0D",
		1709 =>	x"0D0D0D0D",
		1710 =>	x"0D0D0D0D",
		1711 =>	x"0D0D0D0D",
		1712 =>	x"0D0D0D0D",
		1713 =>	x"0D0D0D0D",
		1714 =>	x"0D0D0D0D",
		1715 =>	x"0D0D0D0D",
		1716 =>	x"0D0D0D0D",
		1717 =>	x"0D0D0D0D",
		1718 =>	x"0D0D0D0D",
		1719 =>	x"0D0D0D0D",
		1720 =>	x"0E0E0E0E",
		1721 =>	x"0E0E0E0E",
		1722 =>	x"0E0E0E0E",
		1723 =>	x"0E0E0E0E",
		1724 =>	x"0F0F0F0F",
		1725 =>	x"0F0F0F0F",
		1726 =>	x"0F0F0F0F",
		1727 =>	x"0F0F0F0F",
		1728 =>	x"1011120F", -- IMG_16x16_map_element_18
		1729 =>	x"0F0F0F0F",
		1730 =>	x"0F0F0F0F",
		1731 =>	x"0F121110",
		1732 =>	x"13141516",
		1733 =>	x"0E0E0E0E",
		1734 =>	x"0E0E0E0E",
		1735 =>	x"0E191A11",
		1736 =>	x"12170D0D",
		1737 =>	x"0D0D0D0D",
		1738 =>	x"0D0D0D0D",
		1739 =>	x"0D0D0E12",
		1740 =>	x"0F0E0D0D",
		1741 =>	x"0D0D0D0D",
		1742 =>	x"0D0D0D0D",
		1743 =>	x"0D0D0E0F",
		1744 =>	x"0F0E0D0D",
		1745 =>	x"0D0D0D0D",
		1746 =>	x"0D0D0D0D",
		1747 =>	x"0D0D0E0F",
		1748 =>	x"0F0E0D0D",
		1749 =>	x"0D0D0D0D",
		1750 =>	x"0D0D0D0D",
		1751 =>	x"0D0D0E0F",
		1752 =>	x"0F0E0D0D",
		1753 =>	x"0D0D0D0D",
		1754 =>	x"0D0D0D0D",
		1755 =>	x"0D0D0E0F",
		1756 =>	x"0F0E0D0D",
		1757 =>	x"0D0D0D0D",
		1758 =>	x"0D0D0D0D",
		1759 =>	x"0D0D0E0F",
		1760 =>	x"0F0E0D0D",
		1761 =>	x"0D0D0D0D",
		1762 =>	x"0D0D0D0D",
		1763 =>	x"0D0D0E0F",
		1764 =>	x"0F0E0D0D",
		1765 =>	x"0D0D0D0D",
		1766 =>	x"0D0D0D0D",
		1767 =>	x"0D0D0E0F",
		1768 =>	x"0F0E0D0D",
		1769 =>	x"0D0D0D0D",
		1770 =>	x"0D0D0D0D",
		1771 =>	x"0D0D0E0F",
		1772 =>	x"0F0E0D0D",
		1773 =>	x"0D0D0D0D",
		1774 =>	x"0D0D0D0D",
		1775 =>	x"0D0D0E0F",
		1776 =>	x"0F0E0D0D",
		1777 =>	x"0D0D0D0D",
		1778 =>	x"0D0D0D0D",
		1779 =>	x"0D0D0E0F",
		1780 =>	x"120E0D0D",
		1781 =>	x"0D0D0D0D",
		1782 =>	x"0D0D0D0D",
		1783 =>	x"0D0D0E12",
		1784 =>	x"111A190E",
		1785 =>	x"0E0E0E0E",
		1786 =>	x"0E0E0E0E",
		1787 =>	x"0E191A11",
		1788 =>	x"1011120F",
		1789 =>	x"0F0F0F0F",
		1790 =>	x"0F0F0F0F",
		1791 =>	x"0F121110",
		1792 =>	x"0F0F0F0F", -- IMG_16x16_map_element_19
		1793 =>	x"0F0F0F0F",
		1794 =>	x"0F0F0F0F",
		1795 =>	x"0F0F0F0F",
		1796 =>	x"0E0E0E0E",
		1797 =>	x"0E0E0E0E",
		1798 =>	x"0E0E0E0E",
		1799 =>	x"0E0E0E0E",
		1800 =>	x"0D0D0D0D",
		1801 =>	x"0D0D0D0D",
		1802 =>	x"0D0D0D0D",
		1803 =>	x"0D0D0D0D",
		1804 =>	x"0D0D0D0D",
		1805 =>	x"0D0D0D0D",
		1806 =>	x"0D0D0D0D",
		1807 =>	x"0D0D0D0D",
		1808 =>	x"0D0D0D0D",
		1809 =>	x"0D0D0D0D",
		1810 =>	x"0D0D0D0D",
		1811 =>	x"0D0D0D0D",
		1812 =>	x"0D0D0D0D",
		1813 =>	x"0D0D0D0D",
		1814 =>	x"0D0D0D0D",
		1815 =>	x"0D0D0D0D",
		1816 =>	x"0D0D0D0D",
		1817 =>	x"0D0D0D0D",
		1818 =>	x"0D0D0D0D",
		1819 =>	x"0D0D0D0D",
		1820 =>	x"0D0D0D0D",
		1821 =>	x"0D0D0D0D",
		1822 =>	x"0D0D0D0D",
		1823 =>	x"0D0D0D0D",
		1824 =>	x"0D0D0D0D",
		1825 =>	x"0D0D0D0D",
		1826 =>	x"0D0D0D0D",
		1827 =>	x"0D0D0D0D",
		1828 =>	x"0D0D0D0D",
		1829 =>	x"0D0D0D0D",
		1830 =>	x"0D0D0D0D",
		1831 =>	x"0D0D0D0D",
		1832 =>	x"0D0D0D0D",
		1833 =>	x"0D0D0D0D",
		1834 =>	x"0D0D0D0D",
		1835 =>	x"0D0D0D0D",
		1836 =>	x"0D0D0D0D",
		1837 =>	x"0D0D0D0D",
		1838 =>	x"0D0D0D0D",
		1839 =>	x"0D0D0D0D",
		1840 =>	x"0D0D0D0D",
		1841 =>	x"0D0D0D0D",
		1842 =>	x"0D0D0D0D",
		1843 =>	x"0D0D0D0D",
		1844 =>	x"0D0D0D0D",
		1845 =>	x"0D0D0D0D",
		1846 =>	x"0D0D0D0D",
		1847 =>	x"0D0D0D0D",
		1848 =>	x"0D0D0D0D",
		1849 =>	x"0D0D0D0D",
		1850 =>	x"0D0D0D0D",
		1851 =>	x"0D0D0D0D",
		1852 =>	x"0D0D0D0D",
		1853 =>	x"0D0D0D0D",
		1854 =>	x"0D0D0D0D",
		1855 =>	x"0D0D0D0D",
		1856 =>	x"0F0F0F0F", -- IMG_16x16_map_element_20
		1857 =>	x"0F0F0F0F",
		1858 =>	x"0F0F0F0F",
		1859 =>	x"0F121110",
		1860 =>	x"0E0E0E0E",
		1861 =>	x"0E0E0E0E",
		1862 =>	x"0E0E0E0E",
		1863 =>	x"16151413",
		1864 =>	x"0D0D0D0D",
		1865 =>	x"0D0D0D0D",
		1866 =>	x"0D0D0D0D",
		1867 =>	x"0D0D1712",
		1868 =>	x"0D0D0D0D",
		1869 =>	x"0D0D0D0D",
		1870 =>	x"0D0D0D0D",
		1871 =>	x"0D0D0E0F",
		1872 =>	x"0D0D0D0D",
		1873 =>	x"0D0D0D0D",
		1874 =>	x"0D0D0D0D",
		1875 =>	x"0D0D0E0F",
		1876 =>	x"0D0D0D0D",
		1877 =>	x"0D0D0D0D",
		1878 =>	x"0D0D0D0D",
		1879 =>	x"0D0D0E0F",
		1880 =>	x"0D0D0D0D",
		1881 =>	x"0D0D0D0D",
		1882 =>	x"0D0D0D0D",
		1883 =>	x"0D0D0E0F",
		1884 =>	x"0D0D0D0D",
		1885 =>	x"0D0D0D0D",
		1886 =>	x"0D0D0D0D",
		1887 =>	x"0D0D0E0F",
		1888 =>	x"0D0D0D0D",
		1889 =>	x"0D0D0D0D",
		1890 =>	x"0D0D0D0D",
		1891 =>	x"0D0D0E0F",
		1892 =>	x"0D0D0D0D",
		1893 =>	x"0D0D0D0D",
		1894 =>	x"0D0D0D0D",
		1895 =>	x"0D0D0E0F",
		1896 =>	x"0D0D0D0D",
		1897 =>	x"0D0D0D0D",
		1898 =>	x"0D0D0D0D",
		1899 =>	x"0D0D0E0F",
		1900 =>	x"0D0D0D0D",
		1901 =>	x"0D0D0D0D",
		1902 =>	x"0D0D0D0D",
		1903 =>	x"0D0D0E0F",
		1904 =>	x"0D0D0D0D",
		1905 =>	x"0D0D0D0D",
		1906 =>	x"0D0D0D0D",
		1907 =>	x"0D0D0E0F",
		1908 =>	x"0D0D0D0D",
		1909 =>	x"0D0D0D0D",
		1910 =>	x"0D0D0D0D",
		1911 =>	x"0D0D0E0F",
		1912 =>	x"0D0D0D0D",
		1913 =>	x"0D0D0D0D",
		1914 =>	x"0D0D0D0D",
		1915 =>	x"0D0D0E0F",
		1916 =>	x"0D0D0D0D",
		1917 =>	x"0D0D0D0D",
		1918 =>	x"0D0D0D0D",
		1919 =>	x"0D0D0E0F",
		1920 =>	x"1011120F", -- IMG_16x16_map_element_21
		1921 =>	x"0F0F0F0F",
		1922 =>	x"0F0F0F0F",
		1923 =>	x"0F0F0F0F",
		1924 =>	x"13141516",
		1925 =>	x"0E0E0E0E",
		1926 =>	x"0E0E0E0E",
		1927 =>	x"0E0E0E0E",
		1928 =>	x"12170D0D",
		1929 =>	x"0D0D0D0D",
		1930 =>	x"0D0D0D0D",
		1931 =>	x"0D0D0D0D",
		1932 =>	x"0F0E0D0D",
		1933 =>	x"0D0D0D0D",
		1934 =>	x"0D0D0D0D",
		1935 =>	x"0D0D0D0D",
		1936 =>	x"0F0E0D0D",
		1937 =>	x"0D0D0D0D",
		1938 =>	x"0D0D0D0D",
		1939 =>	x"0D0D0D0D",
		1940 =>	x"0F0E0D0D",
		1941 =>	x"0D0D0D0D",
		1942 =>	x"0D0D0D0D",
		1943 =>	x"0D0D0D0D",
		1944 =>	x"0F0E0D0D",
		1945 =>	x"0D0D0D0D",
		1946 =>	x"0D0D0D0D",
		1947 =>	x"0D0D0D0D",
		1948 =>	x"0F0E0D0D",
		1949 =>	x"0D0D0D0D",
		1950 =>	x"0D0D0D0D",
		1951 =>	x"0D0D0D0D",
		1952 =>	x"0F0E0D0D",
		1953 =>	x"0D0D0D0D",
		1954 =>	x"0D0D0D0D",
		1955 =>	x"0D0D0D0D",
		1956 =>	x"0F0E0D0D",
		1957 =>	x"0D0D0D0D",
		1958 =>	x"0D0D0D0D",
		1959 =>	x"0D0D0D0D",
		1960 =>	x"0F0E0D0D",
		1961 =>	x"0D0D0D0D",
		1962 =>	x"0D0D0D0D",
		1963 =>	x"0D0D0D0D",
		1964 =>	x"0F0E0D0D",
		1965 =>	x"0D0D0D0D",
		1966 =>	x"0D0D0D0D",
		1967 =>	x"0D0D0D0D",
		1968 =>	x"0F0E0D0D",
		1969 =>	x"0D0D0D0D",
		1970 =>	x"0D0D0D0D",
		1971 =>	x"0D0D0D0D",
		1972 =>	x"0F0E0D0D",
		1973 =>	x"0D0D0D0D",
		1974 =>	x"0D0D0D0D",
		1975 =>	x"0D0D0D0D",
		1976 =>	x"0F0E0D0D",
		1977 =>	x"0D0D0D0D",
		1978 =>	x"0D0D0D0D",
		1979 =>	x"0D0D180E",
		1980 =>	x"0F0E0D0D",
		1981 =>	x"0D0D0D0D",
		1982 =>	x"0D0D0D0D",
		1983 =>	x"0D0D0E0F",
		1984 =>	x"1011120F", -- IMG_16x16_map_element_22
		1985 =>	x"0F0F0F0F",
		1986 =>	x"0F0F0F0F",
		1987 =>	x"0F121110",
		1988 =>	x"13141516",
		1989 =>	x"0E0E0E0E",
		1990 =>	x"0E0E0E0E",
		1991 =>	x"16151413",
		1992 =>	x"12170D0D",
		1993 =>	x"0D0D0D0D",
		1994 =>	x"0D0D0D0D",
		1995 =>	x"0D0D1712",
		1996 =>	x"0F0E0D0D",
		1997 =>	x"0D0D0D0D",
		1998 =>	x"0D0D0D0D",
		1999 =>	x"0D0D0E0F",
		2000 =>	x"0F0E0D0D",
		2001 =>	x"0D0D0D0D",
		2002 =>	x"0D0D0D0D",
		2003 =>	x"0D0D0E0F",
		2004 =>	x"0F0E0D0D",
		2005 =>	x"0D0D0D0D",
		2006 =>	x"0D0D0D0D",
		2007 =>	x"0D0D0E0F",
		2008 =>	x"0F0E0D0D",
		2009 =>	x"0D0D0D0D",
		2010 =>	x"0D0D0D0D",
		2011 =>	x"0D0D0E0F",
		2012 =>	x"0F0E0D0D",
		2013 =>	x"0D0D0D0D",
		2014 =>	x"0D0D0D0D",
		2015 =>	x"0D0D0E0F",
		2016 =>	x"0F0E0D0D",
		2017 =>	x"0D0D0D0D",
		2018 =>	x"0D0D0D0D",
		2019 =>	x"0D0D0E0F",
		2020 =>	x"0F0E0D0D",
		2021 =>	x"0D0D0D0D",
		2022 =>	x"0D0D0D0D",
		2023 =>	x"0D0D0E0F",
		2024 =>	x"0F0E0D0D",
		2025 =>	x"0D0D0D0D",
		2026 =>	x"0D0D0D0D",
		2027 =>	x"0D0D0E0F",
		2028 =>	x"0F0E0D0D",
		2029 =>	x"0D0D0D0D",
		2030 =>	x"0D0D0D0D",
		2031 =>	x"0D0D0E0F",
		2032 =>	x"0F0E0D0D",
		2033 =>	x"0D0D0D0D",
		2034 =>	x"0D0D0D0D",
		2035 =>	x"0D0D0E0F",
		2036 =>	x"0F0E0D0D",
		2037 =>	x"0D0D0D0D",
		2038 =>	x"0D0D0D0D",
		2039 =>	x"0D0D0E0F",
		2040 =>	x"0F0E0D0D",
		2041 =>	x"0D0D0D0D",
		2042 =>	x"0D0D0D0D",
		2043 =>	x"0D0D0E0F",
		2044 =>	x"0F0E0D0D",
		2045 =>	x"0D0D0D0D",
		2046 =>	x"0D0D0D0D",
		2047 =>	x"0D0D0E0F",
		2048 =>	x"0F0F0F0F", -- IMG_16x16_map_element_23
		2049 =>	x"0F0F0F0F",
		2050 =>	x"0F0F0F0F",
		2051 =>	x"0F121110",
		2052 =>	x"0E0E0E0E",
		2053 =>	x"0E0E0E0E",
		2054 =>	x"0E0E0E0E",
		2055 =>	x"16151413",
		2056 =>	x"0D0D0D0D",
		2057 =>	x"0D0D0D0D",
		2058 =>	x"0D0D0D0D",
		2059 =>	x"0D0D1712",
		2060 =>	x"0D0D0D0D",
		2061 =>	x"0D0D0D0D",
		2062 =>	x"0D0D0D0D",
		2063 =>	x"0D0D0E0F",
		2064 =>	x"0D0D0D0D",
		2065 =>	x"0D0D0D0D",
		2066 =>	x"0D0D0D0D",
		2067 =>	x"0D0D0E0F",
		2068 =>	x"0D0D0D0D",
		2069 =>	x"0D0D0D0D",
		2070 =>	x"0D0D0D0D",
		2071 =>	x"0D0D0E0F",
		2072 =>	x"0D0D0D0D",
		2073 =>	x"0D0D0D0D",
		2074 =>	x"0D0D0D0D",
		2075 =>	x"0D0D0E0F",
		2076 =>	x"0D0D0D0D",
		2077 =>	x"0D0D0D0D",
		2078 =>	x"0D0D0D0D",
		2079 =>	x"0D0D0E0F",
		2080 =>	x"0D0D0D0D",
		2081 =>	x"0D0D0D0D",
		2082 =>	x"0D0D0D0D",
		2083 =>	x"0D0D0E0F",
		2084 =>	x"0D0D0D0D",
		2085 =>	x"0D0D0D0D",
		2086 =>	x"0D0D0D0D",
		2087 =>	x"0D0D0E0F",
		2088 =>	x"0D0D0D0D",
		2089 =>	x"0D0D0D0D",
		2090 =>	x"0D0D0D0D",
		2091 =>	x"0D0D0E0F",
		2092 =>	x"0D0D0D0D",
		2093 =>	x"0D0D0D0D",
		2094 =>	x"0D0D0D0D",
		2095 =>	x"0D0D0E0F",
		2096 =>	x"0D0D0D0D",
		2097 =>	x"0D0D0D0D",
		2098 =>	x"0D0D0D0D",
		2099 =>	x"0D0D0E0F",
		2100 =>	x"0D0D0D0D",
		2101 =>	x"0D0D0D0D",
		2102 =>	x"0D0D0D0D",
		2103 =>	x"0D0D0E0F",
		2104 =>	x"0E180D0D",
		2105 =>	x"0D0D0D0D",
		2106 =>	x"0D0D0D0D",
		2107 =>	x"0D0D0E0F",
		2108 =>	x"0F0E0D0D",
		2109 =>	x"0D0D0D0D",
		2110 =>	x"0D0D0D0D",
		2111 =>	x"0D0D0E0F",
		2112 =>	x"0F0E0D0D", -- IMG_16x16_map_element_24
		2113 =>	x"0D0D0D0D",
		2114 =>	x"0D0D0D0D",
		2115 =>	x"0D0D0D0D",
		2116 =>	x"0F0E0D0D",
		2117 =>	x"0D0D0D0D",
		2118 =>	x"0D0D0D0D",
		2119 =>	x"0D0D0D0D",
		2120 =>	x"0F0E0D0D",
		2121 =>	x"0D0D0D0D",
		2122 =>	x"0D0D0D0D",
		2123 =>	x"0D0D0D0D",
		2124 =>	x"0F0E0D0D",
		2125 =>	x"0D0D0D0D",
		2126 =>	x"0D0D0D0D",
		2127 =>	x"0D0D0D0D",
		2128 =>	x"0F0E0D0D",
		2129 =>	x"0D0D0D0D",
		2130 =>	x"0D0D0D0D",
		2131 =>	x"0D0D0D0D",
		2132 =>	x"0F0E0D0D",
		2133 =>	x"0D0D0D0D",
		2134 =>	x"0D0D0D0D",
		2135 =>	x"0D0D0D0D",
		2136 =>	x"0F0E0D0D",
		2137 =>	x"0D0D0D0D",
		2138 =>	x"0D0D0D0D",
		2139 =>	x"0D0D0D0D",
		2140 =>	x"0F0E0D0D",
		2141 =>	x"0D0D0D0D",
		2142 =>	x"0D0D0D0D",
		2143 =>	x"0D0D0D0D",
		2144 =>	x"0F0E0D0D",
		2145 =>	x"0D0D0D0D",
		2146 =>	x"0D0D0D0D",
		2147 =>	x"0D0D0D0D",
		2148 =>	x"0F0E0D0D",
		2149 =>	x"0D0D0D0D",
		2150 =>	x"0D0D0D0D",
		2151 =>	x"0D0D0D0D",
		2152 =>	x"0F0E0D0D",
		2153 =>	x"0D0D0D0D",
		2154 =>	x"0D0D0D0D",
		2155 =>	x"0D0D0D0D",
		2156 =>	x"0F0E0D0D",
		2157 =>	x"0D0D0D0D",
		2158 =>	x"0D0D0D0D",
		2159 =>	x"0D0D0D0D",
		2160 =>	x"0F0E0D0D",
		2161 =>	x"0D0D0D0D",
		2162 =>	x"0D0D0D0D",
		2163 =>	x"0D0D0D0D",
		2164 =>	x"0F0E0D0D",
		2165 =>	x"0D0D0D0D",
		2166 =>	x"0D0D0D0D",
		2167 =>	x"0D0D0D0D",
		2168 =>	x"0F0E0D0D",
		2169 =>	x"0D0D0D0D",
		2170 =>	x"0D0D0D0D",
		2171 =>	x"0D0D0D0D",
		2172 =>	x"0F0E0D0D",
		2173 =>	x"0D0D0D0D",
		2174 =>	x"0D0D0D0D",
		2175 =>	x"0D0D0D0D",
		2176 =>	x"0D0D0D0D", -- IMG_16x16_map_element_25
		2177 =>	x"0D0D0D0D",
		2178 =>	x"0D0D0D0D",
		2179 =>	x"0D0D0D0D",
		2180 =>	x"0D0D0D0D",
		2181 =>	x"0D0D0D0D",
		2182 =>	x"0D0D0D0D",
		2183 =>	x"0D0D0D0D",
		2184 =>	x"0D0D0D0D",
		2185 =>	x"0D0D0D0D",
		2186 =>	x"0D0D0D0D",
		2187 =>	x"0D0D0D0D",
		2188 =>	x"0D0D0D0D",
		2189 =>	x"0D0D0D0D",
		2190 =>	x"0D0D0D0D",
		2191 =>	x"0D0D0D0D",
		2192 =>	x"0D0D0D0D",
		2193 =>	x"0D0D0D0D",
		2194 =>	x"0D0D0D0D",
		2195 =>	x"0D0D0D0D",
		2196 =>	x"0D0D0D0D",
		2197 =>	x"0D0D0D0D",
		2198 =>	x"0D0D0D0D",
		2199 =>	x"0D0D0D0D",
		2200 =>	x"0D0D0D0D",
		2201 =>	x"0D0D0D0D",
		2202 =>	x"0D0D0D0D",
		2203 =>	x"0D0D0D0D",
		2204 =>	x"0D0D0D0D",
		2205 =>	x"0D0D0D0D",
		2206 =>	x"0D0D0D0D",
		2207 =>	x"0D0D0D0D",
		2208 =>	x"0D0D0D0D",
		2209 =>	x"0D0D0D0D",
		2210 =>	x"0D0D0D0D",
		2211 =>	x"0D0D0D0D",
		2212 =>	x"0D0D0D0D",
		2213 =>	x"0D0D0D0D",
		2214 =>	x"0D0D0D0D",
		2215 =>	x"0D0D0D0D",
		2216 =>	x"0D0D0D0D",
		2217 =>	x"0D0D0D0D",
		2218 =>	x"0D0D0D0D",
		2219 =>	x"0D0D0D0D",
		2220 =>	x"0D0D0D0D",
		2221 =>	x"0D0D0D0D",
		2222 =>	x"0D0D0D0D",
		2223 =>	x"0D0D0D0D",
		2224 =>	x"0D0D0D0D",
		2225 =>	x"0D0D0D0D",
		2226 =>	x"0D0D0D0D",
		2227 =>	x"0D0D0D0D",
		2228 =>	x"0D0D0D0D",
		2229 =>	x"0D0D0D0D",
		2230 =>	x"0D0D0D0D",
		2231 =>	x"0D0D0D0D",
		2232 =>	x"0D0D0D0D",
		2233 =>	x"0D0D0D0D",
		2234 =>	x"0D0D0D0D",
		2235 =>	x"0D0D0D0D",
		2236 =>	x"0D0D0D0D",
		2237 =>	x"0D0D0D0D",
		2238 =>	x"0D0D0D0D",
		2239 =>	x"0D0D0D0D",
		2240 =>	x"02020202", -- IMG_16x16_rock
		2241 =>	x"02020202",
		2242 =>	x"02020202",
		2243 =>	x"02020202",
		2244 =>	x"02020202",
		2245 =>	x"02000000",
		2246 =>	x"00000202",
		2247 =>	x"02020202",
		2248 =>	x"02020202",
		2249 =>	x"000A0A0A",
		2250 =>	x"0A0A0002",
		2251 =>	x"02020202",
		2252 =>	x"02020200",
		2253 =>	x"0A0A0A0A",
		2254 =>	x"0A0A0002",
		2255 =>	x"02020202",
		2256 =>	x"02020000",
		2257 =>	x"0A0A0A0A",
		2258 =>	x"0A000002",
		2259 =>	x"02020202",
		2260 =>	x"0202000A",
		2261 =>	x"0A000000",
		2262 =>	x"0A0A0A00",
		2263 =>	x"00000002",
		2264 =>	x"0200000A",
		2265 =>	x"0A0A0A00",
		2266 =>	x"0A0A0A0A",
		2267 =>	x"0A0A0000",
		2268 =>	x"000A0000",
		2269 =>	x"00000A00",
		2270 =>	x"0A0A0A00",
		2271 =>	x"0A0A0A00",
		2272 =>	x"000A0A0A",
		2273 =>	x"000A0A00",
		2274 =>	x"0A0A0A0A",
		2275 =>	x"000A0000",
		2276 =>	x"00000A0A",
		2277 =>	x"000A0000",
		2278 =>	x"0A000A0A",
		2279 =>	x"000A0A00",
		2280 =>	x"02000A0A",
		2281 =>	x"000A0A00",
		2282 =>	x"0A0A0A0A",
		2283 =>	x"0A0A0002",
		2284 =>	x"000A0A0A",
		2285 =>	x"000A0A0A",
		2286 =>	x"000A0A00",
		2287 =>	x"00000002",
		2288 =>	x"000A0A0A",
		2289 =>	x"0A0A0A00",
		2290 =>	x"000A0000",
		2291 =>	x"02020202",
		2292 =>	x"0200000A",
		2293 =>	x"0A0A0A00",
		2294 =>	x"0A0A0A00",
		2295 =>	x"02020202",
		2296 =>	x"0202000A",
		2297 =>	x"0A0A0A0A",
		2298 =>	x"0A0A0002",
		2299 =>	x"02020202",
		2300 =>	x"02020200",
		2301 =>	x"0000000A",
		2302 =>	x"00000202",
		2303 =>	x"02020202",
		2304 =>	x"02020202", -- IMG_16x16_smoke
		2305 =>	x"02020202",
		2306 =>	x"02020202",
		2307 =>	x"02020202",
		2308 =>	x"02020200",
		2309 =>	x"00000002",
		2310 =>	x"02020202",
		2311 =>	x"02000002",
		2312 =>	x"02020006",
		2313 =>	x"06060000",
		2314 =>	x"00000002",
		2315 =>	x"00060600",
		2316 =>	x"02000606",
		2317 =>	x"06060006",
		2318 =>	x"06060602",
		2319 =>	x"00060600",
		2320 =>	x"02000006",
		2321 =>	x"06060606",
		2322 =>	x"06060600",
		2323 =>	x"06060600",
		2324 =>	x"06060606",
		2325 =>	x"06000000",
		2326 =>	x"06060000",
		2327 =>	x"06060002",
		2328 =>	x"06060606",
		2329 =>	x"00060606",
		2330 =>	x"00060606",
		2331 =>	x"06060600",
		2332 =>	x"02060600",
		2333 =>	x"06060606",
		2334 =>	x"00000006",
		2335 =>	x"06060600",
		2336 =>	x"06060600",
		2337 =>	x"06060606",
		2338 =>	x"06060006",
		2339 =>	x"06060600",
		2340 =>	x"00060606",
		2341 =>	x"06060606",
		2342 =>	x"06060006",
		2343 =>	x"06060202",
		2344 =>	x"06060606",
		2345 =>	x"06060606",
		2346 =>	x"06060006",
		2347 =>	x"00000002",
		2348 =>	x"02000606",
		2349 =>	x"06060606",
		2350 =>	x"06060006",
		2351 =>	x"06060602",
		2352 =>	x"02000606",
		2353 =>	x"06060606",
		2354 =>	x"00060606",
		2355 =>	x"06060002",
		2356 =>	x"00060606",
		2357 =>	x"06000606",
		2358 =>	x"00060606",
		2359 =>	x"06060002",
		2360 =>	x"00000000",
		2361 =>	x"00000606",
		2362 =>	x"00060606",
		2363 =>	x"06000002",
		2364 =>	x"02020202",
		2365 =>	x"02020000",
		2366 =>	x"02020000",
		2367 =>	x"00020202",


--			***** MAP *****


		2368 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2369 =>	x"00000140", -- z: 0 rot: 0 ptr: 320
		2370 =>	x"00000180", -- z: 0 rot: 0 ptr: 384
		2371 =>	x"000001C0", -- z: 0 rot: 0 ptr: 448
		2372 =>	x"00000200", -- z: 0 rot: 0 ptr: 512
		2373 =>	x"00000240", -- z: 0 rot: 0 ptr: 576
		2374 =>	x"00000280", -- z: 0 rot: 0 ptr: 640
		2375 =>	x"000002C0", -- z: 0 rot: 0 ptr: 704
		2376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2377 =>	x"00000340", -- z: 0 rot: 0 ptr: 832
		2378 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2379 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2380 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2381 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2382 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2383 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2384 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2385 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2386 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2387 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2388 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2389 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2390 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2391 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2392 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2393 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2394 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2395 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2396 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2397 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2398 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2399 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2400 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2401 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2402 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2403 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2404 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2405 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2406 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2407 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2408 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2409 =>	x"00000380", -- z: 0 rot: 0 ptr: 896
		2410 =>	x"000003C0", -- z: 0 rot: 0 ptr: 960
		2411 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2412 =>	x"00000440", -- z: 0 rot: 0 ptr: 1088
		2413 =>	x"00000480", -- z: 0 rot: 0 ptr: 1152
		2414 =>	x"000004C0", -- z: 0 rot: 0 ptr: 1216
		2415 =>	x"00000500", -- z: 0 rot: 0 ptr: 1280
		2416 =>	x"00000540", -- z: 0 rot: 0 ptr: 1344
		2417 =>	x"00000580", -- z: 0 rot: 0 ptr: 1408
		2418 =>	x"000005C0", -- z: 0 rot: 0 ptr: 1472
		2419 =>	x"00000600", -- z: 0 rot: 0 ptr: 1536
		2420 =>	x"00000640", -- z: 0 rot: 0 ptr: 1600
		2421 =>	x"00000680", -- z: 0 rot: 0 ptr: 1664
		2422 =>	x"000006C0", -- z: 0 rot: 0 ptr: 1728
		2423 =>	x"00000700", -- z: 0 rot: 0 ptr: 1792
		2424 =>	x"00000740", -- z: 0 rot: 0 ptr: 1856
		2425 =>	x"000007C0", -- z: 0 rot: 0 ptr: 1984
		2426 =>	x"00000800", -- z: 0 rot: 0 ptr: 2048
		2427 =>	x"00000840", -- z: 0 rot: 0 ptr: 2112
		2428 =>	x"00000880", -- z: 0 rot: 0 ptr: 2176
		2429 =>	x"000004C0", -- z: 0 rot: 0 ptr: 1216
		2430 =>	x"00000600", -- z: 0 rot: 0 ptr: 1536
		2431 =>	x"000008C0", -- z: 0 rot: 0 ptr: 2240
		2432 =>	x"00000900", -- z: 0 rot: 0 ptr: 2304
		2433 =>	x"00000780", -- z: 0 rot: 0 ptr: 1920
		2434 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2435 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2436 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2437 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2438 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2439 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2440 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2441 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2442 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2443 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2444 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2445 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2446 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2447 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2448 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2449 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2450 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2451 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2452 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2453 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2454 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2455 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2456 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2457 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2458 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2459 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2460 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2461 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2462 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2463 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2464 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2465 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2466 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2467 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2468 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2469 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2470 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2471 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2472 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2473 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2474 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2475 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2476 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2477 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2478 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2479 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2480 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2481 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2482 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2483 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2484 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2485 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2486 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2487 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2488 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2489 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2490 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2491 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2492 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2493 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2494 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2495 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2496 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2497 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2498 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2499 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2500 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2501 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2502 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2503 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2504 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2505 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2506 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2507 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2508 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2509 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2510 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2511 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2512 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2513 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2514 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2515 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2516 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2517 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2518 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2519 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2520 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2521 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2522 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2523 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2524 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2525 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2526 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2527 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2528 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2529 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2530 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2531 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2532 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2533 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2534 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2535 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2536 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2537 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2538 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2539 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2540 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2541 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2542 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2543 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2544 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2545 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2546 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2547 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2548 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2549 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2550 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2551 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2552 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2553 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2554 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2555 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2556 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2557 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2558 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2559 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2560 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2561 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2562 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2563 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2564 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2565 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2566 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2567 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2568 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2569 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2570 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2571 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2572 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2573 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2574 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2575 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2576 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2577 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2578 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2579 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2580 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2581 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2582 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2583 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2584 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2585 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2586 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2587 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2588 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2589 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2590 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2591 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2592 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2593 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2594 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2595 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2596 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2597 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2598 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2599 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2600 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2601 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2602 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2603 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2604 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2605 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2606 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2607 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2608 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2609 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2610 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2611 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2612 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2613 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2614 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2615 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2616 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2617 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2618 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2619 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2620 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2621 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2622 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2623 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2624 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2625 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2626 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2627 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2628 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2629 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2630 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2631 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2632 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2633 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2634 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2635 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2636 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2637 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2638 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2639 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2640 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2641 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2642 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2643 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2644 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2645 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2646 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2647 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2648 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2649 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2650 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2651 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2652 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2653 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2654 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2655 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2656 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2657 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2658 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2659 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2660 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2661 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2662 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2663 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2664 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2665 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2666 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2667 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2668 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2669 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2670 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2671 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2672 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2673 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2674 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2675 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2676 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2677 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2678 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2679 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2680 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2681 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2682 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2683 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2684 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2685 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2686 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2687 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2688 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2689 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2690 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2691 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2692 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2693 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2694 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2695 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2696 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2697 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2698 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2699 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2700 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2701 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2702 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2703 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2704 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2705 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2706 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2707 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2708 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2709 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2710 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2711 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2712 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2713 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2714 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2715 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2716 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2717 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2718 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2719 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2720 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2721 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2722 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2723 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2724 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2725 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2726 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2727 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2728 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2729 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2730 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2731 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2732 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2733 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2734 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2735 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2736 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2737 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2738 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2739 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2740 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2741 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2742 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2743 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2744 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2745 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2746 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2747 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2748 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2749 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2750 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2751 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2752 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2753 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2754 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2755 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2756 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2757 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2758 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2759 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2760 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2761 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2762 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2763 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2764 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2765 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2766 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2767 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2768 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2769 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2770 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2771 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2772 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2773 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2774 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2775 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2776 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2777 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2778 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2779 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2780 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2781 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2782 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2783 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2784 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2785 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2786 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2787 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2788 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2789 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2790 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2791 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2792 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2793 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2794 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2795 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2796 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2797 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2798 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2799 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2800 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2801 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2802 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2803 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2804 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2805 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2806 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2807 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2808 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2809 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2810 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2811 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2812 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2813 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2814 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2815 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2816 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2817 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2818 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2819 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2820 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2821 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2822 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2823 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2824 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2825 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2826 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2827 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2828 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2829 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2830 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2831 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2832 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2833 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2834 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2835 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2836 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2837 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2838 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2839 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2840 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2841 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2842 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2843 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2844 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2845 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2846 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2847 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2848 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2849 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2850 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2851 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2852 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2853 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2854 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2855 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2856 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2857 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2858 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2859 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2860 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2861 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2862 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2863 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2864 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2865 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2866 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2867 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2868 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2869 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2870 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2871 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2872 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2873 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2874 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2875 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2876 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2877 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2878 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2879 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2880 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2881 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2882 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2883 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2884 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2885 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2886 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2887 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2888 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2889 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2890 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2891 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2892 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2893 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2894 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2895 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2896 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2897 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2898 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2899 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2900 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2901 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2902 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2903 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2904 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2905 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2906 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2907 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2908 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2909 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2910 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2911 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2912 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2913 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2914 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2915 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2916 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2917 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2918 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2919 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2920 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2921 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2922 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2923 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2924 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2925 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2926 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2927 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2928 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2929 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2930 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2931 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2932 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2933 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2934 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2935 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2936 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2937 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2938 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2939 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2940 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2941 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2942 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2943 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2944 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2945 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2946 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2947 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2948 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2949 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2950 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2951 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2952 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2953 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2954 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2955 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2956 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2957 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2958 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2959 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2960 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2961 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2962 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2963 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2964 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2965 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2966 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2967 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2968 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2969 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2970 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2971 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2972 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2973 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2974 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2975 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2976 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2977 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2978 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2979 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2980 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2981 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2982 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2983 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2984 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2985 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2986 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2987 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2988 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2989 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2990 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2991 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2992 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2993 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2994 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2995 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2996 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2997 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2998 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2999 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3000 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3001 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3002 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3003 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3004 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3005 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3006 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3007 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3008 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3009 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3010 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3011 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3012 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3013 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3014 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3015 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3016 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3017 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3018 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3019 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3020 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3021 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3022 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3023 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3024 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3025 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3026 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3027 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3028 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3029 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3030 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3031 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3032 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3033 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3034 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3035 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3036 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3037 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3038 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3039 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3040 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3041 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3042 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3043 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3044 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3045 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3046 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3047 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3048 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3049 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3050 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3051 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3052 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3053 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3054 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3055 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3056 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3057 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3058 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3059 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3060 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3061 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3062 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3063 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3064 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3065 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3066 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3067 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3068 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3069 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3070 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3071 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3072 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3073 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3074 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3075 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3076 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3077 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3078 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3079 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3080 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3081 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3082 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3083 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3084 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3085 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3086 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3087 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3088 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3089 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3090 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3091 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3092 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3093 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3094 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3095 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3096 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3097 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3098 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3099 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3100 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3101 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3102 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3103 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3104 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3105 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3106 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3107 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3108 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3109 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3110 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3111 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3112 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3113 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3114 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3115 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3116 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3117 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3118 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3119 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3120 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3121 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3122 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3123 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3124 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3125 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3126 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3127 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3128 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3129 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3130 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3131 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3132 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3133 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3134 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3135 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3136 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3137 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3138 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3139 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3140 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3141 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3142 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3143 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3144 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3145 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3146 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3147 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3148 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3149 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3150 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3151 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3152 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3153 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3154 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3155 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3156 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3157 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3158 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3159 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3160 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3161 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3162 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3163 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3164 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3165 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3166 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3167 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3168 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3169 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3170 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3171 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3172 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3173 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3174 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3175 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3176 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3177 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3178 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3179 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3180 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3181 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3182 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3183 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3184 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3185 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3186 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3187 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3188 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3189 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3190 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3191 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3192 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3193 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3194 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3195 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3196 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3197 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3198 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3199 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3200 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3201 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3202 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3203 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3204 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3205 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3206 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3207 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3208 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3209 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3210 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3211 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3212 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3213 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3214 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3215 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3216 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3217 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3218 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3219 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3220 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3221 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3222 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3223 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3224 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3225 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3226 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3227 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3228 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3229 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3230 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3231 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3232 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3233 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3234 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3235 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3236 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3237 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3238 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3239 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3240 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3241 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3242 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3243 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3244 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3245 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3246 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3247 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3248 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3249 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3250 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3251 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3252 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3253 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3254 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3255 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3256 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3257 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3258 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3259 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3260 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3261 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3262 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3263 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3264 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3265 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3266 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3267 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3268 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3269 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3270 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3271 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3272 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3273 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3274 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3275 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3276 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3277 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3278 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3279 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3280 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3281 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3282 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3283 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3284 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3285 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3286 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3287 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3288 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3289 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3290 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3291 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3292 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3293 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3294 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3295 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3296 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3297 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3298 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3299 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3300 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3301 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3302 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3303 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3304 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3305 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3306 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3307 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3308 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3309 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3310 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3311 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3312 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3313 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3314 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3315 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3316 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3317 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3318 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3319 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3320 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3321 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3322 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3323 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3324 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3325 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3326 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3327 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3328 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3329 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3330 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3331 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3332 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3333 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3334 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3335 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3336 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3337 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3338 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3339 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3340 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3341 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3342 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3343 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3344 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3345 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3346 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3347 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3348 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3349 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3350 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3351 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3352 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3353 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3354 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3355 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3356 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3357 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3358 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3359 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3360 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3361 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3362 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3363 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3364 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3365 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3366 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3367 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3368 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3369 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3370 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3371 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3372 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3373 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3374 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3375 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3376 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3377 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3378 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3379 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3380 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3381 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3382 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3383 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3384 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3385 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3386 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3387 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3388 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3389 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3390 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3391 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3392 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3393 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3394 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3395 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3396 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3397 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3398 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3399 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3400 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3401 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3402 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3403 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3404 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3405 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3406 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3407 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3408 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3409 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3410 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3411 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3412 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3413 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3414 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3415 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3416 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3417 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3418 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3419 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3420 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3421 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3422 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3423 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3424 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3425 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3426 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3427 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3428 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3429 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3430 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3431 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3432 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3433 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3434 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3435 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3436 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3437 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3438 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3439 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3440 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3441 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3442 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3443 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3444 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3445 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3446 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3447 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3448 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3449 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3450 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3451 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3452 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3453 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3454 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3455 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3456 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3457 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3458 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3459 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3460 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3461 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3462 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3463 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3464 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3465 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3466 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3467 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3468 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3469 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3470 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3471 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3472 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3473 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3474 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3475 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3476 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3477 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3478 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3479 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3480 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3481 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3482 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3483 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3484 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3485 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3486 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3487 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3488 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3489 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3490 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3491 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3492 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3493 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3494 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3495 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3496 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3497 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3498 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3499 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3500 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3501 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3502 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3503 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3504 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3505 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3506 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3507 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3508 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3509 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3510 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3511 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3512 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3513 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3514 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3515 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3516 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3517 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3518 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3519 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3520 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3521 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3522 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3523 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3524 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3525 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3526 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3527 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3528 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3529 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3530 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3531 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3532 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3533 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3534 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3535 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3536 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3537 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3538 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3539 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3540 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3541 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3542 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3543 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3544 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3545 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3546 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3547 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3548 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3549 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3550 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3551 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3552 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3553 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3554 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3555 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3556 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3557 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3558 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3559 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3560 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3561 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3562 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3563 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3564 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3565 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3566 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3567 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3568 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3569 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3570 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3571 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3572 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3573 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3574 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3575 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3576 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3577 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3578 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3579 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3580 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3581 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3582 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3583 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3584 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3585 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3586 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3587 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3588 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3589 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3590 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3591 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3592 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3593 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3594 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3595 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3596 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3597 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3598 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3599 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3600 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3601 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3602 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3603 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3604 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3605 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3606 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3607 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3608 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3609 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3610 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3611 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3612 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3613 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3614 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3615 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3616 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3617 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3618 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3619 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3620 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3621 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3622 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3623 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3624 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3625 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3626 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3627 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3628 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3629 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3630 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3631 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3632 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3633 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3634 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3635 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3636 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3637 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3638 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		others => x"00000000"
	);

begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;