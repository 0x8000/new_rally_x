
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER
-- DATE: Mon May 14 10:21:16 2018

	signal mem : ram_t := (  -- TODO: Promeniti velicinu mem. Choice 8192 is out of range 0 to 8191 for the index subtype.
	
--			***** COLOR PALLETE *****


		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00277FFF", -- R: 255 G: 127 B: 39
		2 =>	x"0008AF1F", -- R: 31 G: 175 B: 8
		3 =>	x"0000C08F", -- R: 143 G: 192 B: 0
		4 =>	x"001B0080", -- R: 128 G: 0 B: 27
		5 =>	x"00AF1F00", -- R: 0 G: 31 B: 175
		6 =>	x"00E8AF1F", -- R: 31 G: 175 B: 232
		7 =>	x"0000A0AF", -- R: 175 G: 160 B: 0
		8 =>	x"001F0000", -- R: 0 G: 0 B: 31
		9 =>	x"00000070", -- R: 112 G: 0 B: 0
		10 =>	x"00B21F00", -- R: 0 G: 31 B: 178
		11 =>	x"0000AE48", -- R: 72 G: 174 B: 0
		12 =>	x"00B146A8", -- R: 168 G: 70 B: 177
		13 =>	x"00D1000C", -- R: 12 G: 0 B: 209
		14 =>	x"003F0E00", -- R: 0 G: 14 B: 63
		15 =>	x"00000904", -- R: 4 G: 9 B: 0
		16 =>	x"00010000", -- R: 0 G: 0 B: 1
		17 =>	x"00000080", -- R: 128 G: 0 B: 0
		18 =>	x"00AE1F00", -- R: 0 G: 31 B: 174
		19 =>	x"00000600", -- R: 0 G: 6 B: 0
		20 =>	x"000006B8", -- R: 184 G: 6 B: 0
		21 =>	x"00D10000", -- R: 0 G: 0 B: 209
		22 =>	x"0068EF1F", -- R: 31 G: 239 B: 104
		23 =>	x"000060B0", -- R: 176 G: 96 B: 0
		24 =>	x"00530074", -- R: 116 G: 0 B: 83
		25 =>	x"00007500", -- R: 0 G: 117 B: 0
		26 =>	x"00660066", -- R: 102 G: 0 B: 102
		27 =>	x"00005C00", -- R: 0 G: 92 B: 0
		28 =>	x"00310036", -- R: 54 G: 0 B: 49
		29 =>	x"00007800", -- R: 0 G: 120 B: 0
		30 =>	x"003C002E", -- R: 46 G: 0 B: 60
		31 =>	x"00006200", -- R: 0 G: 98 B: 0
		32 =>	x"006D0070", -- R: 112 G: 0 B: 109
		33 =>	x"00B8B31F", -- R: 31 G: 179 B: 184
		34 =>	x"001F0037", -- R: 55 G: 0 B: 31
		35 =>	x"00000037", -- R: 55 G: 0 B: 0
		36 =>	x"00D9D100", -- R: 0 G: 209 B: 217
		37 =>	x"0000B8B3", -- R: 179 G: 184 B: 0
		38 =>	x"001F0060", -- R: 96 G: 0 B: 31
		39 =>	x"00B01F00", -- R: 0 G: 31 B: 176
		40 =>	x"005F006D", -- R: 109 G: 0 B: 95
		41 =>	x"00006500", -- R: 0 G: 101 B: 0
		42 =>	x"006D005C", -- R: 92 G: 0 B: 109
		43 =>	x"00006700", -- R: 0 G: 103 B: 0
		44 =>	x"00720061", -- R: 97 G: 0 B: 114
		45 =>	x"00007000", -- R: 0 G: 112 B: 0
		46 =>	x"00680069", -- R: 105 G: 0 B: 104
		47 =>	x"00006300", -- R: 0 G: 99 B: 0
		48 =>	x"00DDDDDD", -- R: 221 G: 221 B: 221
		49 =>	x"00DD3900", -- R: 0 G: 57 B: 221
		50 =>	x"000039DF", -- R: 223 G: 57 B: 0
		51 =>	x"00FDFDFD", -- R: 253 G: 253 B: 253
		52 =>	x"00FDDDDD", -- R: 221 G: 221 B: 253
		53 =>	x"00DDDDF5", -- R: 245 G: 221 B: 221
		54 =>	x"0048B01C", -- R: 28 G: 176 B: 72
		55 =>	x"00FBD100", -- R: 0 G: 209 B: 251
		56 =>	x"004798FF", -- R: 255 G: 152 B: 71
		57 =>	x"00FF0000", -- R: 0 G: 0 B: 255
		58 =>	x"0000FFFF", -- R: 255 G: 255 B: 0
		59 =>	x"000000FF", -- R: 255 G: 0 B: 0
		60 =>	x"00007F00", -- R: 0 G: 127 B: 0
		61 =>	x"004C4C4C", -- R: 76 G: 76 B: 76
		62 =>	x"007F007F", -- R: 127 G: 0 B: 127
		63 =>	x"0000007F", -- R: 127 G: 0 B: 0
		64 =>	x"00007F82", -- R: 130 G: 127 B: 0
		65 =>	x"00666666", -- R: 102 G: 102 B: 102
		66 =>	x"00DD1F00", -- R: 0 G: 31 B: 221
		67 =>	x"0060B01F", -- R: 31 G: 176 B: 96
		68 =>	x"00003600", -- R: 0 G: 54 B: 0
		69 =>	x"000036D8", -- R: 216 G: 54 B: 0
		70 =>	x"001F005C", -- R: 92 G: 0 B: 31
		71 =>	x"001F00DD", -- R: 221 G: 0 B: 31
		72 =>	x"00000000", -- Unused
		73 =>	x"00000000", -- Unused
		74 =>	x"00000000", -- Unused
		75 =>	x"00000000", -- Unused
		76 =>	x"00000000", -- Unused
		77 =>	x"00000000", -- Unused
		78 =>	x"00000000", -- Unused
		79 =>	x"00000000", -- Unused
		80 =>	x"00000000", -- Unused
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
		255 =>	x"00000000", -- Unused


--			***** 16x16 IMAGES *****


		256 =>	x"01010101", -- IMG_16x16_background
		257 =>	x"01010101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01010101",
		261 =>	x"01010101",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01010101",
		265 =>	x"01010101",
		266 =>	x"01010101",
		267 =>	x"01010101",
		268 =>	x"01010101",
		269 =>	x"01010101",
		270 =>	x"01010101",
		271 =>	x"01010101",
		272 =>	x"01010101",
		273 =>	x"01010101",
		274 =>	x"01010101",
		275 =>	x"01010101",
		276 =>	x"01010101",
		277 =>	x"01010101",
		278 =>	x"01010101",
		279 =>	x"01010101",
		280 =>	x"01010101",
		281 =>	x"01010101",
		282 =>	x"01010101",
		283 =>	x"01010101",
		284 =>	x"01010101",
		285 =>	x"01010101",
		286 =>	x"01010101",
		287 =>	x"01010101",
		288 =>	x"01010101",
		289 =>	x"01010101",
		290 =>	x"01010101",
		291 =>	x"01010101",
		292 =>	x"01010101",
		293 =>	x"01010101",
		294 =>	x"01010101",
		295 =>	x"01010101",
		296 =>	x"01010101",
		297 =>	x"01010101",
		298 =>	x"01010101",
		299 =>	x"01010101",
		300 =>	x"01010101",
		301 =>	x"01010101",
		302 =>	x"01010101",
		303 =>	x"01010101",
		304 =>	x"01010101",
		305 =>	x"01010101",
		306 =>	x"01010101",
		307 =>	x"01010101",
		308 =>	x"01010101",
		309 =>	x"01010101",
		310 =>	x"01010101",
		311 =>	x"01010101",
		312 =>	x"01010101",
		313 =>	x"01010101",
		314 =>	x"01010101",
		315 =>	x"01010101",
		316 =>	x"01010101",
		317 =>	x"01010101",
		318 =>	x"01010101",
		319 =>	x"01010101",
		320 =>	x"02030405", -- IMG_16x16_bang
		321 =>	x"06070800",
		322 =>	x"0000090A",
		323 =>	x"00000000",
		324 =>	x"00000000",
		325 =>	x"000B0C0D",
		326 =>	x"0E0F0000",
		327 =>	x"10001112",
		328 =>	x"00000000",
		329 =>	x"00131415",
		330 =>	x"16170800",
		331 =>	x"00000000",
		332 =>	x"00000000",
		333 =>	x"00000000",
		334 =>	x"00000000",
		335 =>	x"00000000",
		336 =>	x"00000000",
		337 =>	x"00000000",
		338 =>	x"00000000",
		339 =>	x"00000000",
		340 =>	x"00000000",
		341 =>	x"00000000",
		342 =>	x"00000000",
		343 =>	x"00000000",
		344 =>	x"00000000",
		345 =>	x"00000000",
		346 =>	x"00000000",
		347 =>	x"00000000",
		348 =>	x"00000000",
		349 =>	x"00000000",
		350 =>	x"00000000",
		351 =>	x"00000000",
		352 =>	x"00000000",
		353 =>	x"00000000",
		354 =>	x"00000000",
		355 =>	x"00000000",
		356 =>	x"18191A1B",
		357 =>	x"1C1D1C1B",
		358 =>	x"1E1F2000",
		359 =>	x"00000000",
		360 =>	x"21172223",
		361 =>	x"24252627",
		362 =>	x"28292A2B",
		363 =>	x"2C2D2E2F",
		364 =>	x"30303030",
		365 =>	x"30303030",
		366 =>	x"30303030",
		367 =>	x"30313215",
		368 =>	x"30303030",
		369 =>	x"30303030",
		370 =>	x"30303030",
		371 =>	x"30303030",
		372 =>	x"30303030",
		373 =>	x"30303030",
		374 =>	x"30303030",
		375 =>	x"30303030",
		376 =>	x"30303030",
		377 =>	x"30303030",
		378 =>	x"30303030",
		379 =>	x"30303030",
		380 =>	x"33343536",
		381 =>	x"37252627",
		382 =>	x"30303030",
		383 =>	x"30303030",
		384 =>	x"38383838", -- IMG_16x16_car_blue
		385 =>	x"38383838",
		386 =>	x"38383838",
		387 =>	x"38383838",
		388 =>	x"38380000",
		389 =>	x"00383838",
		390 =>	x"38383838",
		391 =>	x"38383838",
		392 =>	x"38380000",
		393 =>	x"00383839",
		394 =>	x"38383838",
		395 =>	x"38383838",
		396 =>	x"38383800",
		397 =>	x"38383839",
		398 =>	x"39383838",
		399 =>	x"38383838",
		400 =>	x"38383939",
		401 =>	x"39393939",
		402 =>	x"39393838",
		403 =>	x"00000038",
		404 =>	x"38000039",
		405 =>	x"39393939",
		406 =>	x"39393939",
		407 =>	x"00000038",
		408 =>	x"38000000",
		409 =>	x"003A3A3A",
		410 =>	x"39393939",
		411 =>	x"38003838",
		412 =>	x"38383939",
		413 =>	x"393A3A3A",
		414 =>	x"3A393939",
		415 =>	x"39393938",
		416 =>	x"38383939",
		417 =>	x"393A3A3A",
		418 =>	x"3A393939",
		419 =>	x"39393938",
		420 =>	x"38000000",
		421 =>	x"003A3A3A",
		422 =>	x"39393939",
		423 =>	x"38003838",
		424 =>	x"38000039",
		425 =>	x"39393939",
		426 =>	x"39393939",
		427 =>	x"00000038",
		428 =>	x"38383939",
		429 =>	x"39393939",
		430 =>	x"39393838",
		431 =>	x"00000038",
		432 =>	x"38383800",
		433 =>	x"38383839",
		434 =>	x"39383838",
		435 =>	x"38383838",
		436 =>	x"38380000",
		437 =>	x"00383839",
		438 =>	x"38383838",
		439 =>	x"38383838",
		440 =>	x"38380000",
		441 =>	x"00383838",
		442 =>	x"38383838",
		443 =>	x"38383838",
		444 =>	x"38383838",
		445 =>	x"38383838",
		446 =>	x"38383838",
		447 =>	x"38383838",
		448 =>	x"38383838", -- IMG_16x16_car_red
		449 =>	x"38383838",
		450 =>	x"38383838",
		451 =>	x"38383838",
		452 =>	x"38380000",
		453 =>	x"00383838",
		454 =>	x"38383838",
		455 =>	x"38383838",
		456 =>	x"38380000",
		457 =>	x"0038383B",
		458 =>	x"38383838",
		459 =>	x"38383838",
		460 =>	x"38383800",
		461 =>	x"3838383B",
		462 =>	x"3B383838",
		463 =>	x"38383838",
		464 =>	x"38383B3B",
		465 =>	x"3B3B3B3B",
		466 =>	x"3B3B3838",
		467 =>	x"00000038",
		468 =>	x"3800003B",
		469 =>	x"3B3B3B3B",
		470 =>	x"3B3B3B3B",
		471 =>	x"00000038",
		472 =>	x"38000000",
		473 =>	x"003A3A3A",
		474 =>	x"3B3B3B3B",
		475 =>	x"38003838",
		476 =>	x"38383B3B",
		477 =>	x"3B3A3A3A",
		478 =>	x"3A3B3B3B",
		479 =>	x"3B3B3B38",
		480 =>	x"38383B3B",
		481 =>	x"3B3A3A3A",
		482 =>	x"3A3B3B3B",
		483 =>	x"3B3B3B38",
		484 =>	x"38000000",
		485 =>	x"003A3A3A",
		486 =>	x"3B3B3B3B",
		487 =>	x"38003838",
		488 =>	x"3800003B",
		489 =>	x"3B3B3B3B",
		490 =>	x"3B3B3B3B",
		491 =>	x"00000038",
		492 =>	x"38383B3B",
		493 =>	x"3B3B3B3B",
		494 =>	x"3B3B3838",
		495 =>	x"00000038",
		496 =>	x"38383800",
		497 =>	x"3838383B",
		498 =>	x"3B383838",
		499 =>	x"38383838",
		500 =>	x"38380000",
		501 =>	x"0038383B",
		502 =>	x"38383838",
		503 =>	x"38383838",
		504 =>	x"38380000",
		505 =>	x"00383838",
		506 =>	x"38383838",
		507 =>	x"38383838",
		508 =>	x"38383838",
		509 =>	x"38383838",
		510 =>	x"38383838",
		511 =>	x"38383838",
		512 =>	x"01010101", -- IMG_16x16_flag
		513 =>	x"01010101",
		514 =>	x"01010101",
		515 =>	x"01010101",
		516 =>	x"01013A3A",
		517 =>	x"01010101",
		518 =>	x"01010101",
		519 =>	x"01010101",
		520 =>	x"01013A3A",
		521 =>	x"3A3A0101",
		522 =>	x"01010101",
		523 =>	x"01010101",
		524 =>	x"01013A3A",
		525 =>	x"3A3A3A3A",
		526 =>	x"01010101",
		527 =>	x"01010101",
		528 =>	x"01013A3A",
		529 =>	x"3A3A3A3A",
		530 =>	x"3A3A0101",
		531 =>	x"01010101",
		532 =>	x"01013A3A",
		533 =>	x"3A3A3A3A",
		534 =>	x"3A3A3A3A",
		535 =>	x"01010101",
		536 =>	x"01013A3A",
		537 =>	x"3A3A3A3A",
		538 =>	x"3A3A0101",
		539 =>	x"01010101",
		540 =>	x"01013A3A",
		541 =>	x"3A3A3A3A",
		542 =>	x"01010101",
		543 =>	x"01010101",
		544 =>	x"01013A3A",
		545 =>	x"3A3A0101",
		546 =>	x"01010101",
		547 =>	x"01010101",
		548 =>	x"01013A3A",
		549 =>	x"01010101",
		550 =>	x"01010101",
		551 =>	x"01010101",
		552 =>	x"01013A3A",
		553 =>	x"01010101",
		554 =>	x"01010101",
		555 =>	x"01010101",
		556 =>	x"01013A3A",
		557 =>	x"01010101",
		558 =>	x"01010101",
		559 =>	x"01010101",
		560 =>	x"01013A3A",
		561 =>	x"01010101",
		562 =>	x"01010101",
		563 =>	x"01010101",
		564 =>	x"013A3A3A",
		565 =>	x"3A010101",
		566 =>	x"01010101",
		567 =>	x"01010101",
		568 =>	x"013A3A3A",
		569 =>	x"3A010101",
		570 =>	x"01010101",
		571 =>	x"01010101",
		572 =>	x"01010101",
		573 =>	x"01010101",
		574 =>	x"01010101",
		575 =>	x"01010101",
		576 =>	x"3C3C3C3C", -- IMG_16x16_map_element_00
		577 =>	x"3C3C3D3C",
		578 =>	x"3D3D3C3C",
		579 =>	x"3C3C3C3C",
		580 =>	x"3C3C3C3C",
		581 =>	x"3E3F3F3E",
		582 =>	x"3F3E3F3D",
		583 =>	x"3C3C3C3C",
		584 =>	x"3C3C3D3F",
		585 =>	x"3E3F3F3E",
		586 =>	x"40413F3F",
		587 =>	x"3C3C3C3C",
		588 =>	x"3C3C3E3F",
		589 =>	x"3F3F3E3E",
		590 =>	x"3F3F3E3E",
		591 =>	x"3F3F3C3C",
		592 =>	x"3C3D3F3F",
		593 =>	x"3F3F3E3E",
		594 =>	x"3F3B3E3E",
		595 =>	x"3E3D3D3C",
		596 =>	x"3D3E3E3F",
		597 =>	x"3F3B3E3E",
		598 =>	x"3F3B3E3F",
		599 =>	x"3F3F3F3D",
		600 =>	x"3D3F3F3F",
		601 =>	x"3F3F3F3E",
		602 =>	x"3F3F3F3B",
		603 =>	x"3B3F3F3D",
		604 =>	x"3D403E3E",
		605 =>	x"3F3E3E3D",
		606 =>	x"3E3E3F3E",
		607 =>	x"3B3F3D3D",
		608 =>	x"3D3F3F40",
		609 =>	x"3F3F3F3F",
		610 =>	x"3F3F3F3B",
		611 =>	x"3F3F3F3D",
		612 =>	x"3D3F3F3F",
		613 =>	x"3F403F3E",
		614 =>	x"3F3F3E3F",
		615 =>	x"3E3F3E3D",
		616 =>	x"3D3E3F3F",
		617 =>	x"3F3F3E3F",
		618 =>	x"3B3E3F3F",
		619 =>	x"3E3D3E3D",
		620 =>	x"3C3F3F3E",
		621 =>	x"3E3E3E3F",
		622 =>	x"3F3E3E3F",
		623 =>	x"3E3E3D3C",
		624 =>	x"3C3C3E3F",
		625 =>	x"3F3E3F3F",
		626 =>	x"3E3E3E3F",
		627 =>	x"3F3F3D3C",
		628 =>	x"3C3C3D40",
		629 =>	x"3F3E403F",
		630 =>	x"3E3E3F3F",
		631 =>	x"3E3D3C3C",
		632 =>	x"3C3C3C3C",
		633 =>	x"3D3F4040",
		634 =>	x"3F3B3D3C",
		635 =>	x"3C3C3C3C",
		636 =>	x"3C3C3C3C",
		637 =>	x"3C3C3D3D",
		638 =>	x"3D3D3C3C",
		639 =>	x"3C3C3C3C",
		640 =>	x"02030405", -- IMG_16x16_map_element_01
		641 =>	x"06070800",
		642 =>	x"0000090A",
		643 =>	x"00000000",
		644 =>	x"00000000",
		645 =>	x"000B0C0D",
		646 =>	x"0E0F0000",
		647 =>	x"10001112",
		648 =>	x"00000000",
		649 =>	x"00131415",
		650 =>	x"16170800",
		651 =>	x"00000000",
		652 =>	x"00000000",
		653 =>	x"00000000",
		654 =>	x"00000000",
		655 =>	x"00000000",
		656 =>	x"00000000",
		657 =>	x"00000000",
		658 =>	x"00000000",
		659 =>	x"00000000",
		660 =>	x"00000000",
		661 =>	x"00000000",
		662 =>	x"00000000",
		663 =>	x"00000000",
		664 =>	x"00000000",
		665 =>	x"00000000",
		666 =>	x"00000000",
		667 =>	x"00000000",
		668 =>	x"00000000",
		669 =>	x"00000000",
		670 =>	x"00000000",
		671 =>	x"00000000",
		672 =>	x"00000000",
		673 =>	x"00000000",
		674 =>	x"00000000",
		675 =>	x"00000000",
		676 =>	x"18191A1B",
		677 =>	x"1C1D1C1B",
		678 =>	x"1E1F2000",
		679 =>	x"00000000",
		680 =>	x"30303042",
		681 =>	x"43444515",
		682 =>	x"2117462B",
		683 =>	x"2C2D2E2F",
		684 =>	x"30303030",
		685 =>	x"30303030",
		686 =>	x"30303030",
		687 =>	x"30303030",
		688 =>	x"30303030",
		689 =>	x"30303030",
		690 =>	x"30303030",
		691 =>	x"30303030",
		692 =>	x"30303030",
		693 =>	x"30303030",
		694 =>	x"30303030",
		695 =>	x"30303030",
		696 =>	x"30303030",
		697 =>	x"30303030",
		698 =>	x"30303030",
		699 =>	x"30303030",
		700 =>	x"33343536",
		701 =>	x"37252627",
		702 =>	x"30303030",
		703 =>	x"30303030",
		704 =>	x"02030405", -- IMG_16x16_map_element_02
		705 =>	x"06070800",
		706 =>	x"0000090A",
		707 =>	x"00000000",
		708 =>	x"00000000",
		709 =>	x"000B0C0D",
		710 =>	x"0E0F0000",
		711 =>	x"10001112",
		712 =>	x"00000000",
		713 =>	x"00131415",
		714 =>	x"16170800",
		715 =>	x"00000000",
		716 =>	x"00000000",
		717 =>	x"00000000",
		718 =>	x"00000000",
		719 =>	x"00000000",
		720 =>	x"00000000",
		721 =>	x"00000000",
		722 =>	x"00000000",
		723 =>	x"00000000",
		724 =>	x"00000000",
		725 =>	x"00000000",
		726 =>	x"00000000",
		727 =>	x"00000000",
		728 =>	x"00000000",
		729 =>	x"00000000",
		730 =>	x"00000000",
		731 =>	x"00000000",
		732 =>	x"00000000",
		733 =>	x"00000000",
		734 =>	x"00000000",
		735 =>	x"00000000",
		736 =>	x"00000000",
		737 =>	x"00000000",
		738 =>	x"00000000",
		739 =>	x"00000000",
		740 =>	x"18191A1B",
		741 =>	x"1C1D1C1B",
		742 =>	x"1E1F2000",
		743 =>	x"00000000",
		744 =>	x"30303042",
		745 =>	x"43444515",
		746 =>	x"2117462B",
		747 =>	x"2C2D2E2F",
		748 =>	x"30303030",
		749 =>	x"30303030",
		750 =>	x"30303030",
		751 =>	x"30303030",
		752 =>	x"30303030",
		753 =>	x"30303030",
		754 =>	x"30303030",
		755 =>	x"30303030",
		756 =>	x"30303030",
		757 =>	x"30303030",
		758 =>	x"30303030",
		759 =>	x"30303030",
		760 =>	x"30303030",
		761 =>	x"30303030",
		762 =>	x"30303030",
		763 =>	x"30303030",
		764 =>	x"33343536",
		765 =>	x"37252627",
		766 =>	x"30303030",
		767 =>	x"30303030",
		768 =>	x"02030405", -- IMG_16x16_map_element_03
		769 =>	x"06070800",
		770 =>	x"0000090A",
		771 =>	x"00000000",
		772 =>	x"00000000",
		773 =>	x"000B0C0D",
		774 =>	x"0E0F0000",
		775 =>	x"10001112",
		776 =>	x"00000000",
		777 =>	x"00131415",
		778 =>	x"16170800",
		779 =>	x"00000000",
		780 =>	x"00000000",
		781 =>	x"00000000",
		782 =>	x"00000000",
		783 =>	x"00000000",
		784 =>	x"00000000",
		785 =>	x"00000000",
		786 =>	x"00000000",
		787 =>	x"00000000",
		788 =>	x"00000000",
		789 =>	x"00000000",
		790 =>	x"00000000",
		791 =>	x"00000000",
		792 =>	x"00000000",
		793 =>	x"00000000",
		794 =>	x"00000000",
		795 =>	x"00000000",
		796 =>	x"00000000",
		797 =>	x"00000000",
		798 =>	x"00000000",
		799 =>	x"00000000",
		800 =>	x"00000000",
		801 =>	x"00000000",
		802 =>	x"00000000",
		803 =>	x"00000000",
		804 =>	x"18191A1B",
		805 =>	x"1C1D1C1B",
		806 =>	x"1E1F2000",
		807 =>	x"00000000",
		808 =>	x"30303042",
		809 =>	x"43444515",
		810 =>	x"2117462B",
		811 =>	x"2C2D2E2F",
		812 =>	x"30303030",
		813 =>	x"30303030",
		814 =>	x"30303030",
		815 =>	x"30303030",
		816 =>	x"30303030",
		817 =>	x"30303030",
		818 =>	x"30303030",
		819 =>	x"30303030",
		820 =>	x"30303030",
		821 =>	x"30303030",
		822 =>	x"30303030",
		823 =>	x"30303030",
		824 =>	x"30303030",
		825 =>	x"30303030",
		826 =>	x"30303030",
		827 =>	x"30303030",
		828 =>	x"33343536",
		829 =>	x"37252627",
		830 =>	x"30303030",
		831 =>	x"30303030",
		832 =>	x"02030405", -- IMG_16x16_map_element_04
		833 =>	x"06070800",
		834 =>	x"0000090A",
		835 =>	x"00000000",
		836 =>	x"00000000",
		837 =>	x"000B0C0D",
		838 =>	x"0E0F0000",
		839 =>	x"10001112",
		840 =>	x"00000000",
		841 =>	x"00131415",
		842 =>	x"16170800",
		843 =>	x"00000000",
		844 =>	x"00000000",
		845 =>	x"00000000",
		846 =>	x"00000000",
		847 =>	x"00000000",
		848 =>	x"00000000",
		849 =>	x"00000000",
		850 =>	x"00000000",
		851 =>	x"00000000",
		852 =>	x"00000000",
		853 =>	x"00000000",
		854 =>	x"00000000",
		855 =>	x"00000000",
		856 =>	x"00000000",
		857 =>	x"00000000",
		858 =>	x"00000000",
		859 =>	x"00000000",
		860 =>	x"00000000",
		861 =>	x"00000000",
		862 =>	x"00000000",
		863 =>	x"00000000",
		864 =>	x"00000000",
		865 =>	x"00000000",
		866 =>	x"00000000",
		867 =>	x"00000000",
		868 =>	x"18191A1B",
		869 =>	x"1C1D1C1B",
		870 =>	x"1E1F2000",
		871 =>	x"00000000",
		872 =>	x"30303042",
		873 =>	x"43444515",
		874 =>	x"2117462B",
		875 =>	x"2C2D2E2F",
		876 =>	x"30303030",
		877 =>	x"30303030",
		878 =>	x"30303030",
		879 =>	x"30303030",
		880 =>	x"30303030",
		881 =>	x"30303030",
		882 =>	x"30303030",
		883 =>	x"30303030",
		884 =>	x"30303030",
		885 =>	x"30303030",
		886 =>	x"30303030",
		887 =>	x"30303030",
		888 =>	x"30303030",
		889 =>	x"30303030",
		890 =>	x"30303030",
		891 =>	x"30303030",
		892 =>	x"33343536",
		893 =>	x"37252627",
		894 =>	x"30303030",
		895 =>	x"30303030",
		896 =>	x"02030405", -- IMG_16x16_map_element_05
		897 =>	x"06070800",
		898 =>	x"0000090A",
		899 =>	x"00000000",
		900 =>	x"00000000",
		901 =>	x"000B0C0D",
		902 =>	x"0E0F0000",
		903 =>	x"10001112",
		904 =>	x"00000000",
		905 =>	x"00131415",
		906 =>	x"16170800",
		907 =>	x"00000000",
		908 =>	x"00000000",
		909 =>	x"00000000",
		910 =>	x"00000000",
		911 =>	x"00000000",
		912 =>	x"00000000",
		913 =>	x"00000000",
		914 =>	x"00000000",
		915 =>	x"00000000",
		916 =>	x"00000000",
		917 =>	x"00000000",
		918 =>	x"00000000",
		919 =>	x"00000000",
		920 =>	x"00000000",
		921 =>	x"00000000",
		922 =>	x"00000000",
		923 =>	x"00000000",
		924 =>	x"00000000",
		925 =>	x"00000000",
		926 =>	x"00000000",
		927 =>	x"00000000",
		928 =>	x"00000000",
		929 =>	x"00000000",
		930 =>	x"00000000",
		931 =>	x"00000000",
		932 =>	x"18191A1B",
		933 =>	x"1C1D1C1B",
		934 =>	x"1E1F2000",
		935 =>	x"00000000",
		936 =>	x"30303042",
		937 =>	x"43444515",
		938 =>	x"2117462B",
		939 =>	x"2C2D2E2F",
		940 =>	x"30303030",
		941 =>	x"30303030",
		942 =>	x"30303030",
		943 =>	x"30303030",
		944 =>	x"30303030",
		945 =>	x"30303030",
		946 =>	x"30303030",
		947 =>	x"30303030",
		948 =>	x"30303030",
		949 =>	x"30303030",
		950 =>	x"30303030",
		951 =>	x"30303030",
		952 =>	x"30303030",
		953 =>	x"30303030",
		954 =>	x"30303030",
		955 =>	x"30303030",
		956 =>	x"33343536",
		957 =>	x"37252627",
		958 =>	x"30303030",
		959 =>	x"30303030",
		960 =>	x"02030405", -- IMG_16x16_map_element_06
		961 =>	x"06070800",
		962 =>	x"0000090A",
		963 =>	x"00000000",
		964 =>	x"00000000",
		965 =>	x"000B0C0D",
		966 =>	x"0E0F0000",
		967 =>	x"10001112",
		968 =>	x"00000000",
		969 =>	x"00131415",
		970 =>	x"16170800",
		971 =>	x"00000000",
		972 =>	x"00000000",
		973 =>	x"00000000",
		974 =>	x"00000000",
		975 =>	x"00000000",
		976 =>	x"00000000",
		977 =>	x"00000000",
		978 =>	x"00000000",
		979 =>	x"00000000",
		980 =>	x"00000000",
		981 =>	x"00000000",
		982 =>	x"00000000",
		983 =>	x"00000000",
		984 =>	x"00000000",
		985 =>	x"00000000",
		986 =>	x"00000000",
		987 =>	x"00000000",
		988 =>	x"00000000",
		989 =>	x"00000000",
		990 =>	x"00000000",
		991 =>	x"00000000",
		992 =>	x"00000000",
		993 =>	x"00000000",
		994 =>	x"00000000",
		995 =>	x"00000000",
		996 =>	x"18191A1B",
		997 =>	x"1C1D1C1B",
		998 =>	x"1E1F2000",
		999 =>	x"00000000",
		1000 =>	x"30303042",
		1001 =>	x"43444515",
		1002 =>	x"2117462B",
		1003 =>	x"2C2D2E2F",
		1004 =>	x"30303030",
		1005 =>	x"30303030",
		1006 =>	x"30303030",
		1007 =>	x"30303030",
		1008 =>	x"30303030",
		1009 =>	x"30303030",
		1010 =>	x"30303030",
		1011 =>	x"30303030",
		1012 =>	x"30303030",
		1013 =>	x"30303030",
		1014 =>	x"30303030",
		1015 =>	x"30303030",
		1016 =>	x"30303030",
		1017 =>	x"30303030",
		1018 =>	x"30303030",
		1019 =>	x"30303030",
		1020 =>	x"33343536",
		1021 =>	x"37252627",
		1022 =>	x"30303030",
		1023 =>	x"30303030",
		1024 =>	x"02030405", -- IMG_16x16_map_element_07
		1025 =>	x"06070800",
		1026 =>	x"0000090A",
		1027 =>	x"00000000",
		1028 =>	x"00000000",
		1029 =>	x"000B0C0D",
		1030 =>	x"0E0F0000",
		1031 =>	x"10001112",
		1032 =>	x"00000000",
		1033 =>	x"00131415",
		1034 =>	x"16170800",
		1035 =>	x"00000000",
		1036 =>	x"00000000",
		1037 =>	x"00000000",
		1038 =>	x"00000000",
		1039 =>	x"00000000",
		1040 =>	x"00000000",
		1041 =>	x"00000000",
		1042 =>	x"00000000",
		1043 =>	x"00000000",
		1044 =>	x"00000000",
		1045 =>	x"00000000",
		1046 =>	x"00000000",
		1047 =>	x"00000000",
		1048 =>	x"00000000",
		1049 =>	x"00000000",
		1050 =>	x"00000000",
		1051 =>	x"00000000",
		1052 =>	x"00000000",
		1053 =>	x"00000000",
		1054 =>	x"00000000",
		1055 =>	x"00000000",
		1056 =>	x"00000000",
		1057 =>	x"00000000",
		1058 =>	x"00000000",
		1059 =>	x"00000000",
		1060 =>	x"18191A1B",
		1061 =>	x"1C1D1C1B",
		1062 =>	x"1E1F2000",
		1063 =>	x"00000000",
		1064 =>	x"30303042",
		1065 =>	x"43444515",
		1066 =>	x"2117462B",
		1067 =>	x"2C2D2E2F",
		1068 =>	x"30303030",
		1069 =>	x"30303030",
		1070 =>	x"30303030",
		1071 =>	x"30303030",
		1072 =>	x"30303030",
		1073 =>	x"30303030",
		1074 =>	x"30303030",
		1075 =>	x"30303030",
		1076 =>	x"30303030",
		1077 =>	x"30303030",
		1078 =>	x"30303030",
		1079 =>	x"30303030",
		1080 =>	x"30303030",
		1081 =>	x"30303030",
		1082 =>	x"30303030",
		1083 =>	x"30303030",
		1084 =>	x"33343536",
		1085 =>	x"37252627",
		1086 =>	x"30303030",
		1087 =>	x"30303030",
		1088 =>	x"02030405", -- IMG_16x16_map_element_08
		1089 =>	x"06070800",
		1090 =>	x"0000090A",
		1091 =>	x"00000000",
		1092 =>	x"00000000",
		1093 =>	x"000B0C0D",
		1094 =>	x"0E0F0000",
		1095 =>	x"10001112",
		1096 =>	x"00000000",
		1097 =>	x"00131415",
		1098 =>	x"16170800",
		1099 =>	x"00000000",
		1100 =>	x"00000000",
		1101 =>	x"00000000",
		1102 =>	x"00000000",
		1103 =>	x"00000000",
		1104 =>	x"00000000",
		1105 =>	x"00000000",
		1106 =>	x"00000000",
		1107 =>	x"00000000",
		1108 =>	x"00000000",
		1109 =>	x"00000000",
		1110 =>	x"00000000",
		1111 =>	x"00000000",
		1112 =>	x"00000000",
		1113 =>	x"00000000",
		1114 =>	x"00000000",
		1115 =>	x"00000000",
		1116 =>	x"00000000",
		1117 =>	x"00000000",
		1118 =>	x"00000000",
		1119 =>	x"00000000",
		1120 =>	x"00000000",
		1121 =>	x"00000000",
		1122 =>	x"00000000",
		1123 =>	x"00000000",
		1124 =>	x"18191A1B",
		1125 =>	x"1C1D1C1B",
		1126 =>	x"1E1F2000",
		1127 =>	x"00000000",
		1128 =>	x"30303042",
		1129 =>	x"43444515",
		1130 =>	x"2117462B",
		1131 =>	x"2C2D2E2F",
		1132 =>	x"30303030",
		1133 =>	x"30303030",
		1134 =>	x"30303030",
		1135 =>	x"30303030",
		1136 =>	x"30303030",
		1137 =>	x"30303030",
		1138 =>	x"30303030",
		1139 =>	x"30303030",
		1140 =>	x"30303030",
		1141 =>	x"30303030",
		1142 =>	x"30303030",
		1143 =>	x"30303030",
		1144 =>	x"30303030",
		1145 =>	x"30303030",
		1146 =>	x"30303030",
		1147 =>	x"30303030",
		1148 =>	x"33343536",
		1149 =>	x"37252627",
		1150 =>	x"30303030",
		1151 =>	x"30303030",
		1152 =>	x"02030405", -- IMG_16x16_map_element_09
		1153 =>	x"06070800",
		1154 =>	x"0000090A",
		1155 =>	x"00000000",
		1156 =>	x"00000000",
		1157 =>	x"000B0C0D",
		1158 =>	x"0E0F0000",
		1159 =>	x"10001112",
		1160 =>	x"00000000",
		1161 =>	x"00131415",
		1162 =>	x"16170800",
		1163 =>	x"00000000",
		1164 =>	x"00000000",
		1165 =>	x"00000000",
		1166 =>	x"00000000",
		1167 =>	x"00000000",
		1168 =>	x"00000000",
		1169 =>	x"00000000",
		1170 =>	x"00000000",
		1171 =>	x"00000000",
		1172 =>	x"00000000",
		1173 =>	x"00000000",
		1174 =>	x"00000000",
		1175 =>	x"00000000",
		1176 =>	x"00000000",
		1177 =>	x"00000000",
		1178 =>	x"00000000",
		1179 =>	x"00000000",
		1180 =>	x"00000000",
		1181 =>	x"00000000",
		1182 =>	x"00000000",
		1183 =>	x"00000000",
		1184 =>	x"00000000",
		1185 =>	x"00000000",
		1186 =>	x"00000000",
		1187 =>	x"00000000",
		1188 =>	x"18191A1B",
		1189 =>	x"1C1D1C1B",
		1190 =>	x"1E1F2000",
		1191 =>	x"00000000",
		1192 =>	x"30303042",
		1193 =>	x"43444515",
		1194 =>	x"2117462B",
		1195 =>	x"2C2D2E2F",
		1196 =>	x"30303030",
		1197 =>	x"30303030",
		1198 =>	x"30303030",
		1199 =>	x"30303030",
		1200 =>	x"30303030",
		1201 =>	x"30303030",
		1202 =>	x"30303030",
		1203 =>	x"30303030",
		1204 =>	x"30303030",
		1205 =>	x"30303030",
		1206 =>	x"30303030",
		1207 =>	x"30303030",
		1208 =>	x"30303030",
		1209 =>	x"30303030",
		1210 =>	x"30303030",
		1211 =>	x"30303030",
		1212 =>	x"33343536",
		1213 =>	x"37252627",
		1214 =>	x"30303030",
		1215 =>	x"30303030",
		1216 =>	x"02030405", -- IMG_16x16_map_element_10
		1217 =>	x"06070800",
		1218 =>	x"0000090A",
		1219 =>	x"00000000",
		1220 =>	x"00000000",
		1221 =>	x"000B0C0D",
		1222 =>	x"0E0F0000",
		1223 =>	x"10001112",
		1224 =>	x"00000000",
		1225 =>	x"00131415",
		1226 =>	x"16170800",
		1227 =>	x"00000000",
		1228 =>	x"00000000",
		1229 =>	x"00000000",
		1230 =>	x"00000000",
		1231 =>	x"00000000",
		1232 =>	x"00000000",
		1233 =>	x"00000000",
		1234 =>	x"00000000",
		1235 =>	x"00000000",
		1236 =>	x"00000000",
		1237 =>	x"00000000",
		1238 =>	x"00000000",
		1239 =>	x"00000000",
		1240 =>	x"00000000",
		1241 =>	x"00000000",
		1242 =>	x"00000000",
		1243 =>	x"00000000",
		1244 =>	x"00000000",
		1245 =>	x"00000000",
		1246 =>	x"00000000",
		1247 =>	x"00000000",
		1248 =>	x"00000000",
		1249 =>	x"00000000",
		1250 =>	x"00000000",
		1251 =>	x"00000000",
		1252 =>	x"18191A1B",
		1253 =>	x"1C1D1C1B",
		1254 =>	x"1E1F2000",
		1255 =>	x"00000000",
		1256 =>	x"30303042",
		1257 =>	x"43444515",
		1258 =>	x"2117462B",
		1259 =>	x"2C2D2E2F",
		1260 =>	x"30303030",
		1261 =>	x"30303030",
		1262 =>	x"30303030",
		1263 =>	x"30303030",
		1264 =>	x"30303030",
		1265 =>	x"30303030",
		1266 =>	x"30303030",
		1267 =>	x"30303030",
		1268 =>	x"30303030",
		1269 =>	x"30303030",
		1270 =>	x"30303030",
		1271 =>	x"30303030",
		1272 =>	x"30303030",
		1273 =>	x"30303030",
		1274 =>	x"30303030",
		1275 =>	x"30303030",
		1276 =>	x"33343536",
		1277 =>	x"37252627",
		1278 =>	x"30303030",
		1279 =>	x"30303030",
		1280 =>	x"02030405", -- IMG_16x16_map_element_11
		1281 =>	x"06070800",
		1282 =>	x"0000090A",
		1283 =>	x"00000000",
		1284 =>	x"00000000",
		1285 =>	x"000B0C0D",
		1286 =>	x"0E0F0000",
		1287 =>	x"10001112",
		1288 =>	x"00000000",
		1289 =>	x"00131415",
		1290 =>	x"16170800",
		1291 =>	x"00000000",
		1292 =>	x"00000000",
		1293 =>	x"00000000",
		1294 =>	x"00000000",
		1295 =>	x"00000000",
		1296 =>	x"00000000",
		1297 =>	x"00000000",
		1298 =>	x"00000000",
		1299 =>	x"00000000",
		1300 =>	x"00000000",
		1301 =>	x"00000000",
		1302 =>	x"00000000",
		1303 =>	x"00000000",
		1304 =>	x"00000000",
		1305 =>	x"00000000",
		1306 =>	x"00000000",
		1307 =>	x"00000000",
		1308 =>	x"00000000",
		1309 =>	x"00000000",
		1310 =>	x"00000000",
		1311 =>	x"00000000",
		1312 =>	x"00000000",
		1313 =>	x"00000000",
		1314 =>	x"00000000",
		1315 =>	x"00000000",
		1316 =>	x"18191A1B",
		1317 =>	x"1C1D1C1B",
		1318 =>	x"1E1F2000",
		1319 =>	x"00000000",
		1320 =>	x"30303042",
		1321 =>	x"43444515",
		1322 =>	x"2117462B",
		1323 =>	x"2C2D2E2F",
		1324 =>	x"30303030",
		1325 =>	x"30303030",
		1326 =>	x"30303030",
		1327 =>	x"30303030",
		1328 =>	x"30303030",
		1329 =>	x"30303030",
		1330 =>	x"30303030",
		1331 =>	x"30303030",
		1332 =>	x"30303030",
		1333 =>	x"30303030",
		1334 =>	x"30303030",
		1335 =>	x"30303030",
		1336 =>	x"30303030",
		1337 =>	x"30303030",
		1338 =>	x"30303030",
		1339 =>	x"30303030",
		1340 =>	x"33343536",
		1341 =>	x"37252627",
		1342 =>	x"30303030",
		1343 =>	x"30303030",
		1344 =>	x"02030405", -- IMG_16x16_map_element_12
		1345 =>	x"06070800",
		1346 =>	x"0000090A",
		1347 =>	x"00000000",
		1348 =>	x"00000000",
		1349 =>	x"000B0C0D",
		1350 =>	x"0E0F0000",
		1351 =>	x"10001112",
		1352 =>	x"00000000",
		1353 =>	x"00131415",
		1354 =>	x"16170800",
		1355 =>	x"00000000",
		1356 =>	x"00000000",
		1357 =>	x"00000000",
		1358 =>	x"00000000",
		1359 =>	x"00000000",
		1360 =>	x"00000000",
		1361 =>	x"00000000",
		1362 =>	x"00000000",
		1363 =>	x"00000000",
		1364 =>	x"00000000",
		1365 =>	x"00000000",
		1366 =>	x"00000000",
		1367 =>	x"00000000",
		1368 =>	x"00000000",
		1369 =>	x"00000000",
		1370 =>	x"00000000",
		1371 =>	x"00000000",
		1372 =>	x"00000000",
		1373 =>	x"00000000",
		1374 =>	x"00000000",
		1375 =>	x"00000000",
		1376 =>	x"00000000",
		1377 =>	x"00000000",
		1378 =>	x"00000000",
		1379 =>	x"00000000",
		1380 =>	x"18191A1B",
		1381 =>	x"1C1D1C1B",
		1382 =>	x"1E1F2000",
		1383 =>	x"00000000",
		1384 =>	x"30303042",
		1385 =>	x"43444515",
		1386 =>	x"2117462B",
		1387 =>	x"2C2D2E2F",
		1388 =>	x"30303030",
		1389 =>	x"30303030",
		1390 =>	x"30303030",
		1391 =>	x"30303030",
		1392 =>	x"30303030",
		1393 =>	x"30303030",
		1394 =>	x"30303030",
		1395 =>	x"30303030",
		1396 =>	x"30303030",
		1397 =>	x"30303030",
		1398 =>	x"30303030",
		1399 =>	x"30303030",
		1400 =>	x"30303030",
		1401 =>	x"30303030",
		1402 =>	x"30303030",
		1403 =>	x"30303030",
		1404 =>	x"33343536",
		1405 =>	x"37252627",
		1406 =>	x"30303030",
		1407 =>	x"30303030",
		1408 =>	x"02030405", -- IMG_16x16_map_element_13
		1409 =>	x"06070800",
		1410 =>	x"0000090A",
		1411 =>	x"00000000",
		1412 =>	x"00000000",
		1413 =>	x"000B0C0D",
		1414 =>	x"0E0F0000",
		1415 =>	x"10001112",
		1416 =>	x"00000000",
		1417 =>	x"00131415",
		1418 =>	x"16170800",
		1419 =>	x"00000000",
		1420 =>	x"00000000",
		1421 =>	x"00000000",
		1422 =>	x"00000000",
		1423 =>	x"00000000",
		1424 =>	x"00000000",
		1425 =>	x"00000000",
		1426 =>	x"00000000",
		1427 =>	x"00000000",
		1428 =>	x"00000000",
		1429 =>	x"00000000",
		1430 =>	x"00000000",
		1431 =>	x"00000000",
		1432 =>	x"00000000",
		1433 =>	x"00000000",
		1434 =>	x"00000000",
		1435 =>	x"00000000",
		1436 =>	x"00000000",
		1437 =>	x"00000000",
		1438 =>	x"00000000",
		1439 =>	x"00000000",
		1440 =>	x"00000000",
		1441 =>	x"00000000",
		1442 =>	x"00000000",
		1443 =>	x"00000000",
		1444 =>	x"18191A1B",
		1445 =>	x"1C1D1C1B",
		1446 =>	x"1E1F2000",
		1447 =>	x"00000000",
		1448 =>	x"30303042",
		1449 =>	x"43444515",
		1450 =>	x"2117462B",
		1451 =>	x"2C2D2E2F",
		1452 =>	x"30303030",
		1453 =>	x"30303030",
		1454 =>	x"30303030",
		1455 =>	x"30303030",
		1456 =>	x"30303030",
		1457 =>	x"30303030",
		1458 =>	x"30303030",
		1459 =>	x"30303030",
		1460 =>	x"30303030",
		1461 =>	x"30303030",
		1462 =>	x"30303030",
		1463 =>	x"30303030",
		1464 =>	x"30303030",
		1465 =>	x"30303030",
		1466 =>	x"30303030",
		1467 =>	x"30303030",
		1468 =>	x"33343536",
		1469 =>	x"37252627",
		1470 =>	x"30303030",
		1471 =>	x"30303030",
		1472 =>	x"02030405", -- IMG_16x16_map_element_14
		1473 =>	x"06070800",
		1474 =>	x"0000090A",
		1475 =>	x"00000000",
		1476 =>	x"00000000",
		1477 =>	x"000B0C0D",
		1478 =>	x"0E0F0000",
		1479 =>	x"10001112",
		1480 =>	x"00000000",
		1481 =>	x"00131415",
		1482 =>	x"16170800",
		1483 =>	x"00000000",
		1484 =>	x"00000000",
		1485 =>	x"00000000",
		1486 =>	x"00000000",
		1487 =>	x"00000000",
		1488 =>	x"00000000",
		1489 =>	x"00000000",
		1490 =>	x"00000000",
		1491 =>	x"00000000",
		1492 =>	x"00000000",
		1493 =>	x"00000000",
		1494 =>	x"00000000",
		1495 =>	x"00000000",
		1496 =>	x"00000000",
		1497 =>	x"00000000",
		1498 =>	x"00000000",
		1499 =>	x"00000000",
		1500 =>	x"00000000",
		1501 =>	x"00000000",
		1502 =>	x"00000000",
		1503 =>	x"00000000",
		1504 =>	x"00000000",
		1505 =>	x"00000000",
		1506 =>	x"00000000",
		1507 =>	x"00000000",
		1508 =>	x"18191A1B",
		1509 =>	x"1C1D1C1B",
		1510 =>	x"1E1F2000",
		1511 =>	x"00000000",
		1512 =>	x"30303042",
		1513 =>	x"43444515",
		1514 =>	x"2117462B",
		1515 =>	x"2C2D2E2F",
		1516 =>	x"30303030",
		1517 =>	x"30303030",
		1518 =>	x"30303030",
		1519 =>	x"30303030",
		1520 =>	x"30303030",
		1521 =>	x"30303030",
		1522 =>	x"30303030",
		1523 =>	x"30303030",
		1524 =>	x"30303030",
		1525 =>	x"30303030",
		1526 =>	x"30303030",
		1527 =>	x"30303030",
		1528 =>	x"30303030",
		1529 =>	x"30303030",
		1530 =>	x"30303030",
		1531 =>	x"30303030",
		1532 =>	x"33343536",
		1533 =>	x"37252627",
		1534 =>	x"30303030",
		1535 =>	x"30303030",
		1536 =>	x"02030405", -- IMG_16x16_map_element_15
		1537 =>	x"06070800",
		1538 =>	x"0000090A",
		1539 =>	x"00000000",
		1540 =>	x"00000000",
		1541 =>	x"000B0C0D",
		1542 =>	x"0E0F0000",
		1543 =>	x"10001112",
		1544 =>	x"00000000",
		1545 =>	x"00131415",
		1546 =>	x"16170800",
		1547 =>	x"00000000",
		1548 =>	x"00000000",
		1549 =>	x"00000000",
		1550 =>	x"00000000",
		1551 =>	x"00000000",
		1552 =>	x"00000000",
		1553 =>	x"00000000",
		1554 =>	x"00000000",
		1555 =>	x"00000000",
		1556 =>	x"00000000",
		1557 =>	x"00000000",
		1558 =>	x"00000000",
		1559 =>	x"00000000",
		1560 =>	x"00000000",
		1561 =>	x"00000000",
		1562 =>	x"00000000",
		1563 =>	x"00000000",
		1564 =>	x"00000000",
		1565 =>	x"00000000",
		1566 =>	x"00000000",
		1567 =>	x"00000000",
		1568 =>	x"00000000",
		1569 =>	x"00000000",
		1570 =>	x"00000000",
		1571 =>	x"00000000",
		1572 =>	x"18191A1B",
		1573 =>	x"1C1D1C1B",
		1574 =>	x"1E1F2000",
		1575 =>	x"00000000",
		1576 =>	x"30303042",
		1577 =>	x"43444515",
		1578 =>	x"2117462B",
		1579 =>	x"2C2D2E2F",
		1580 =>	x"30303030",
		1581 =>	x"30303030",
		1582 =>	x"30303030",
		1583 =>	x"30303030",
		1584 =>	x"30303030",
		1585 =>	x"30303030",
		1586 =>	x"30303030",
		1587 =>	x"30303030",
		1588 =>	x"30303030",
		1589 =>	x"30303030",
		1590 =>	x"30303030",
		1591 =>	x"30303030",
		1592 =>	x"30303030",
		1593 =>	x"30303030",
		1594 =>	x"30303030",
		1595 =>	x"30303030",
		1596 =>	x"33343536",
		1597 =>	x"37252627",
		1598 =>	x"30303030",
		1599 =>	x"30303030",
		1600 =>	x"02030405", -- IMG_16x16_map_element_16
		1601 =>	x"06070800",
		1602 =>	x"0000090A",
		1603 =>	x"00000000",
		1604 =>	x"00000000",
		1605 =>	x"000B0C0D",
		1606 =>	x"0E0F0000",
		1607 =>	x"10001112",
		1608 =>	x"00000000",
		1609 =>	x"00131415",
		1610 =>	x"16170800",
		1611 =>	x"00000000",
		1612 =>	x"00000000",
		1613 =>	x"00000000",
		1614 =>	x"00000000",
		1615 =>	x"00000000",
		1616 =>	x"00000000",
		1617 =>	x"00000000",
		1618 =>	x"00000000",
		1619 =>	x"00000000",
		1620 =>	x"00000000",
		1621 =>	x"00000000",
		1622 =>	x"00000000",
		1623 =>	x"00000000",
		1624 =>	x"00000000",
		1625 =>	x"00000000",
		1626 =>	x"00000000",
		1627 =>	x"00000000",
		1628 =>	x"00000000",
		1629 =>	x"00000000",
		1630 =>	x"00000000",
		1631 =>	x"00000000",
		1632 =>	x"00000000",
		1633 =>	x"00000000",
		1634 =>	x"00000000",
		1635 =>	x"00000000",
		1636 =>	x"18191A1B",
		1637 =>	x"1C1D1C1B",
		1638 =>	x"1E1F2000",
		1639 =>	x"00000000",
		1640 =>	x"30303042",
		1641 =>	x"43444515",
		1642 =>	x"2117462B",
		1643 =>	x"2C2D2E2F",
		1644 =>	x"30303030",
		1645 =>	x"30303030",
		1646 =>	x"30303030",
		1647 =>	x"30303030",
		1648 =>	x"30303030",
		1649 =>	x"30303030",
		1650 =>	x"30303030",
		1651 =>	x"30303030",
		1652 =>	x"30303030",
		1653 =>	x"30303030",
		1654 =>	x"30303030",
		1655 =>	x"30303030",
		1656 =>	x"30303030",
		1657 =>	x"30303030",
		1658 =>	x"30303030",
		1659 =>	x"30303030",
		1660 =>	x"33343536",
		1661 =>	x"37252627",
		1662 =>	x"30303030",
		1663 =>	x"30303030",
		1664 =>	x"02030405", -- IMG_16x16_map_element_17
		1665 =>	x"06070800",
		1666 =>	x"0000090A",
		1667 =>	x"00000000",
		1668 =>	x"00000000",
		1669 =>	x"000B0C0D",
		1670 =>	x"0E0F0000",
		1671 =>	x"10001112",
		1672 =>	x"00000000",
		1673 =>	x"00131415",
		1674 =>	x"16170800",
		1675 =>	x"00000000",
		1676 =>	x"00000000",
		1677 =>	x"00000000",
		1678 =>	x"00000000",
		1679 =>	x"00000000",
		1680 =>	x"00000000",
		1681 =>	x"00000000",
		1682 =>	x"00000000",
		1683 =>	x"00000000",
		1684 =>	x"00000000",
		1685 =>	x"00000000",
		1686 =>	x"00000000",
		1687 =>	x"00000000",
		1688 =>	x"00000000",
		1689 =>	x"00000000",
		1690 =>	x"00000000",
		1691 =>	x"00000000",
		1692 =>	x"00000000",
		1693 =>	x"00000000",
		1694 =>	x"00000000",
		1695 =>	x"00000000",
		1696 =>	x"00000000",
		1697 =>	x"00000000",
		1698 =>	x"00000000",
		1699 =>	x"00000000",
		1700 =>	x"18191A1B",
		1701 =>	x"1C1D1C1B",
		1702 =>	x"1E1F2000",
		1703 =>	x"00000000",
		1704 =>	x"30303042",
		1705 =>	x"43444515",
		1706 =>	x"2117462B",
		1707 =>	x"2C2D2E2F",
		1708 =>	x"30303030",
		1709 =>	x"30303030",
		1710 =>	x"30303030",
		1711 =>	x"30303030",
		1712 =>	x"30303030",
		1713 =>	x"30303030",
		1714 =>	x"30303030",
		1715 =>	x"30303030",
		1716 =>	x"30303030",
		1717 =>	x"30303030",
		1718 =>	x"30303030",
		1719 =>	x"30303030",
		1720 =>	x"30303030",
		1721 =>	x"30303030",
		1722 =>	x"30303030",
		1723 =>	x"30303030",
		1724 =>	x"33343536",
		1725 =>	x"37252627",
		1726 =>	x"30303030",
		1727 =>	x"30303030",
		1728 =>	x"02030405", -- IMG_16x16_map_element_18
		1729 =>	x"06070800",
		1730 =>	x"0000090A",
		1731 =>	x"00000000",
		1732 =>	x"00000000",
		1733 =>	x"000B0C0D",
		1734 =>	x"0E0F0000",
		1735 =>	x"10001112",
		1736 =>	x"00000000",
		1737 =>	x"00131415",
		1738 =>	x"16170800",
		1739 =>	x"00000000",
		1740 =>	x"00000000",
		1741 =>	x"00000000",
		1742 =>	x"00000000",
		1743 =>	x"00000000",
		1744 =>	x"00000000",
		1745 =>	x"00000000",
		1746 =>	x"00000000",
		1747 =>	x"00000000",
		1748 =>	x"00000000",
		1749 =>	x"00000000",
		1750 =>	x"00000000",
		1751 =>	x"00000000",
		1752 =>	x"00000000",
		1753 =>	x"00000000",
		1754 =>	x"00000000",
		1755 =>	x"00000000",
		1756 =>	x"00000000",
		1757 =>	x"00000000",
		1758 =>	x"00000000",
		1759 =>	x"00000000",
		1760 =>	x"00000000",
		1761 =>	x"00000000",
		1762 =>	x"00000000",
		1763 =>	x"00000000",
		1764 =>	x"18191A1B",
		1765 =>	x"1C1D1C1B",
		1766 =>	x"1E1F2000",
		1767 =>	x"00000000",
		1768 =>	x"30303042",
		1769 =>	x"43444515",
		1770 =>	x"2117462B",
		1771 =>	x"2C2D2E2F",
		1772 =>	x"30303030",
		1773 =>	x"30303030",
		1774 =>	x"30303030",
		1775 =>	x"30303030",
		1776 =>	x"30303030",
		1777 =>	x"30303030",
		1778 =>	x"30303030",
		1779 =>	x"30303030",
		1780 =>	x"30303030",
		1781 =>	x"30303030",
		1782 =>	x"30303030",
		1783 =>	x"30303030",
		1784 =>	x"30303030",
		1785 =>	x"30303030",
		1786 =>	x"30303030",
		1787 =>	x"30303030",
		1788 =>	x"33343536",
		1789 =>	x"37252627",
		1790 =>	x"30303030",
		1791 =>	x"30303030",
		1792 =>	x"02030405", -- IMG_16x16_map_element_19
		1793 =>	x"06070800",
		1794 =>	x"0000090A",
		1795 =>	x"00000000",
		1796 =>	x"00000000",
		1797 =>	x"000B0C0D",
		1798 =>	x"0E0F0000",
		1799 =>	x"10001112",
		1800 =>	x"00000000",
		1801 =>	x"00131415",
		1802 =>	x"16170800",
		1803 =>	x"00000000",
		1804 =>	x"00000000",
		1805 =>	x"00000000",
		1806 =>	x"00000000",
		1807 =>	x"00000000",
		1808 =>	x"00000000",
		1809 =>	x"00000000",
		1810 =>	x"00000000",
		1811 =>	x"00000000",
		1812 =>	x"00000000",
		1813 =>	x"00000000",
		1814 =>	x"00000000",
		1815 =>	x"00000000",
		1816 =>	x"00000000",
		1817 =>	x"00000000",
		1818 =>	x"00000000",
		1819 =>	x"00000000",
		1820 =>	x"00000000",
		1821 =>	x"00000000",
		1822 =>	x"00000000",
		1823 =>	x"00000000",
		1824 =>	x"00000000",
		1825 =>	x"00000000",
		1826 =>	x"00000000",
		1827 =>	x"00000000",
		1828 =>	x"18191A1B",
		1829 =>	x"1C1D1C1B",
		1830 =>	x"1E1F2000",
		1831 =>	x"00000000",
		1832 =>	x"30303042",
		1833 =>	x"43444515",
		1834 =>	x"2117462B",
		1835 =>	x"2C2D2E2F",
		1836 =>	x"30303030",
		1837 =>	x"30303030",
		1838 =>	x"30303030",
		1839 =>	x"30303030",
		1840 =>	x"30303030",
		1841 =>	x"30303030",
		1842 =>	x"30303030",
		1843 =>	x"30303030",
		1844 =>	x"30303030",
		1845 =>	x"30303030",
		1846 =>	x"30303030",
		1847 =>	x"30303030",
		1848 =>	x"30303030",
		1849 =>	x"30303030",
		1850 =>	x"30303030",
		1851 =>	x"30303030",
		1852 =>	x"33343536",
		1853 =>	x"37252627",
		1854 =>	x"30303030",
		1855 =>	x"30303030",
		1856 =>	x"02030405", -- IMG_16x16_map_element_20
		1857 =>	x"06070800",
		1858 =>	x"0000090A",
		1859 =>	x"00000000",
		1860 =>	x"00000000",
		1861 =>	x"000B0C0D",
		1862 =>	x"0E0F0000",
		1863 =>	x"10001112",
		1864 =>	x"00000000",
		1865 =>	x"00131415",
		1866 =>	x"16170800",
		1867 =>	x"00000000",
		1868 =>	x"00000000",
		1869 =>	x"00000000",
		1870 =>	x"00000000",
		1871 =>	x"00000000",
		1872 =>	x"00000000",
		1873 =>	x"00000000",
		1874 =>	x"00000000",
		1875 =>	x"00000000",
		1876 =>	x"00000000",
		1877 =>	x"00000000",
		1878 =>	x"00000000",
		1879 =>	x"00000000",
		1880 =>	x"00000000",
		1881 =>	x"00000000",
		1882 =>	x"00000000",
		1883 =>	x"00000000",
		1884 =>	x"00000000",
		1885 =>	x"00000000",
		1886 =>	x"00000000",
		1887 =>	x"00000000",
		1888 =>	x"00000000",
		1889 =>	x"00000000",
		1890 =>	x"00000000",
		1891 =>	x"00000000",
		1892 =>	x"18191A1B",
		1893 =>	x"1C1D1C1B",
		1894 =>	x"1E1F2000",
		1895 =>	x"00000000",
		1896 =>	x"30303042",
		1897 =>	x"43444515",
		1898 =>	x"2117462B",
		1899 =>	x"2C2D2E2F",
		1900 =>	x"30303030",
		1901 =>	x"30303030",
		1902 =>	x"30303030",
		1903 =>	x"30303030",
		1904 =>	x"30303030",
		1905 =>	x"30303030",
		1906 =>	x"30303030",
		1907 =>	x"30303030",
		1908 =>	x"30303030",
		1909 =>	x"30303030",
		1910 =>	x"30303030",
		1911 =>	x"30303030",
		1912 =>	x"30303030",
		1913 =>	x"30303030",
		1914 =>	x"30303030",
		1915 =>	x"30303030",
		1916 =>	x"33343536",
		1917 =>	x"37252627",
		1918 =>	x"30303030",
		1919 =>	x"30303030",
		1920 =>	x"02030405", -- IMG_16x16_map_element_21
		1921 =>	x"06070800",
		1922 =>	x"0000090A",
		1923 =>	x"00000000",
		1924 =>	x"00000000",
		1925 =>	x"000B0C0D",
		1926 =>	x"0E0F0000",
		1927 =>	x"10001112",
		1928 =>	x"00000000",
		1929 =>	x"00131415",
		1930 =>	x"16170800",
		1931 =>	x"00000000",
		1932 =>	x"00000000",
		1933 =>	x"00000000",
		1934 =>	x"00000000",
		1935 =>	x"00000000",
		1936 =>	x"00000000",
		1937 =>	x"00000000",
		1938 =>	x"00000000",
		1939 =>	x"00000000",
		1940 =>	x"00000000",
		1941 =>	x"00000000",
		1942 =>	x"00000000",
		1943 =>	x"00000000",
		1944 =>	x"00000000",
		1945 =>	x"00000000",
		1946 =>	x"00000000",
		1947 =>	x"00000000",
		1948 =>	x"00000000",
		1949 =>	x"00000000",
		1950 =>	x"00000000",
		1951 =>	x"00000000",
		1952 =>	x"00000000",
		1953 =>	x"00000000",
		1954 =>	x"00000000",
		1955 =>	x"00000000",
		1956 =>	x"18191A1B",
		1957 =>	x"1C1D1C1B",
		1958 =>	x"1E1F2000",
		1959 =>	x"00000000",
		1960 =>	x"30303042",
		1961 =>	x"43444515",
		1962 =>	x"2117462B",
		1963 =>	x"2C2D2E2F",
		1964 =>	x"30303030",
		1965 =>	x"30303030",
		1966 =>	x"30303030",
		1967 =>	x"30303030",
		1968 =>	x"30303030",
		1969 =>	x"30303030",
		1970 =>	x"30303030",
		1971 =>	x"30303030",
		1972 =>	x"30303030",
		1973 =>	x"30303030",
		1974 =>	x"30303030",
		1975 =>	x"30303030",
		1976 =>	x"30303030",
		1977 =>	x"30303030",
		1978 =>	x"30303030",
		1979 =>	x"30303030",
		1980 =>	x"33343536",
		1981 =>	x"37252627",
		1982 =>	x"30303030",
		1983 =>	x"30303030",
		1984 =>	x"02030405", -- IMG_16x16_map_element_22
		1985 =>	x"06070800",
		1986 =>	x"0000090A",
		1987 =>	x"00000000",
		1988 =>	x"00000000",
		1989 =>	x"000B0C0D",
		1990 =>	x"0E0F0000",
		1991 =>	x"10001112",
		1992 =>	x"00000000",
		1993 =>	x"00131415",
		1994 =>	x"16170800",
		1995 =>	x"00000000",
		1996 =>	x"00000000",
		1997 =>	x"00000000",
		1998 =>	x"00000000",
		1999 =>	x"00000000",
		2000 =>	x"00000000",
		2001 =>	x"00000000",
		2002 =>	x"00000000",
		2003 =>	x"00000000",
		2004 =>	x"00000000",
		2005 =>	x"00000000",
		2006 =>	x"00000000",
		2007 =>	x"00000000",
		2008 =>	x"00000000",
		2009 =>	x"00000000",
		2010 =>	x"00000000",
		2011 =>	x"00000000",
		2012 =>	x"00000000",
		2013 =>	x"00000000",
		2014 =>	x"00000000",
		2015 =>	x"00000000",
		2016 =>	x"00000000",
		2017 =>	x"00000000",
		2018 =>	x"00000000",
		2019 =>	x"00000000",
		2020 =>	x"18191A1B",
		2021 =>	x"1C1D1C1B",
		2022 =>	x"1E1F2000",
		2023 =>	x"00000000",
		2024 =>	x"30303042",
		2025 =>	x"43444515",
		2026 =>	x"2117462B",
		2027 =>	x"2C2D2E2F",
		2028 =>	x"30303030",
		2029 =>	x"30303030",
		2030 =>	x"30303030",
		2031 =>	x"30303030",
		2032 =>	x"30303030",
		2033 =>	x"30303030",
		2034 =>	x"30303030",
		2035 =>	x"30303030",
		2036 =>	x"30303030",
		2037 =>	x"30303030",
		2038 =>	x"30303030",
		2039 =>	x"30303030",
		2040 =>	x"30303030",
		2041 =>	x"30303030",
		2042 =>	x"30303030",
		2043 =>	x"30303030",
		2044 =>	x"33343536",
		2045 =>	x"37252627",
		2046 =>	x"30303030",
		2047 =>	x"30303030",
		2048 =>	x"02030405", -- IMG_16x16_map_element_23
		2049 =>	x"06070800",
		2050 =>	x"0000090A",
		2051 =>	x"00000000",
		2052 =>	x"00000000",
		2053 =>	x"000B0C0D",
		2054 =>	x"0E0F0000",
		2055 =>	x"10001112",
		2056 =>	x"00000000",
		2057 =>	x"00131415",
		2058 =>	x"16170800",
		2059 =>	x"00000000",
		2060 =>	x"00000000",
		2061 =>	x"00000000",
		2062 =>	x"00000000",
		2063 =>	x"00000000",
		2064 =>	x"00000000",
		2065 =>	x"00000000",
		2066 =>	x"00000000",
		2067 =>	x"00000000",
		2068 =>	x"00000000",
		2069 =>	x"00000000",
		2070 =>	x"00000000",
		2071 =>	x"00000000",
		2072 =>	x"00000000",
		2073 =>	x"00000000",
		2074 =>	x"00000000",
		2075 =>	x"00000000",
		2076 =>	x"00000000",
		2077 =>	x"00000000",
		2078 =>	x"00000000",
		2079 =>	x"00000000",
		2080 =>	x"00000000",
		2081 =>	x"00000000",
		2082 =>	x"00000000",
		2083 =>	x"00000000",
		2084 =>	x"18191A1B",
		2085 =>	x"1C1D1C1B",
		2086 =>	x"1E1F2000",
		2087 =>	x"00000000",
		2088 =>	x"30303042",
		2089 =>	x"43444515",
		2090 =>	x"2117462B",
		2091 =>	x"2C2D2E2F",
		2092 =>	x"30303030",
		2093 =>	x"30303030",
		2094 =>	x"30303030",
		2095 =>	x"30303030",
		2096 =>	x"30303030",
		2097 =>	x"30303030",
		2098 =>	x"30303030",
		2099 =>	x"30303030",
		2100 =>	x"30303030",
		2101 =>	x"30303030",
		2102 =>	x"30303030",
		2103 =>	x"30303030",
		2104 =>	x"30303030",
		2105 =>	x"30303030",
		2106 =>	x"30303030",
		2107 =>	x"30303030",
		2108 =>	x"33343536",
		2109 =>	x"37252627",
		2110 =>	x"30303030",
		2111 =>	x"30303030",
		2112 =>	x"02030405", -- IMG_16x16_map_element_24
		2113 =>	x"06070800",
		2114 =>	x"0000090A",
		2115 =>	x"00000000",
		2116 =>	x"00000000",
		2117 =>	x"000B0C0D",
		2118 =>	x"0E0F0000",
		2119 =>	x"10001112",
		2120 =>	x"00000000",
		2121 =>	x"00131415",
		2122 =>	x"16170800",
		2123 =>	x"00000000",
		2124 =>	x"00000000",
		2125 =>	x"00000000",
		2126 =>	x"00000000",
		2127 =>	x"00000000",
		2128 =>	x"00000000",
		2129 =>	x"00000000",
		2130 =>	x"00000000",
		2131 =>	x"00000000",
		2132 =>	x"00000000",
		2133 =>	x"00000000",
		2134 =>	x"00000000",
		2135 =>	x"00000000",
		2136 =>	x"00000000",
		2137 =>	x"00000000",
		2138 =>	x"00000000",
		2139 =>	x"00000000",
		2140 =>	x"00000000",
		2141 =>	x"00000000",
		2142 =>	x"00000000",
		2143 =>	x"00000000",
		2144 =>	x"00000000",
		2145 =>	x"00000000",
		2146 =>	x"00000000",
		2147 =>	x"00000000",
		2148 =>	x"18191A1B",
		2149 =>	x"1C1D1C1B",
		2150 =>	x"1E1F2000",
		2151 =>	x"00000000",
		2152 =>	x"30303042",
		2153 =>	x"43444515",
		2154 =>	x"2117462B",
		2155 =>	x"2C2D2E2F",
		2156 =>	x"30303030",
		2157 =>	x"30303030",
		2158 =>	x"30303030",
		2159 =>	x"30303030",
		2160 =>	x"30303030",
		2161 =>	x"30303030",
		2162 =>	x"30303030",
		2163 =>	x"30303030",
		2164 =>	x"30303030",
		2165 =>	x"30303030",
		2166 =>	x"30303030",
		2167 =>	x"30303030",
		2168 =>	x"30303030",
		2169 =>	x"30303030",
		2170 =>	x"30303030",
		2171 =>	x"30303030",
		2172 =>	x"33343536",
		2173 =>	x"37252627",
		2174 =>	x"30303030",
		2175 =>	x"30303030",
		2176 =>	x"02030405", -- IMG_16x16_map_element_25
		2177 =>	x"06070800",
		2178 =>	x"0000090A",
		2179 =>	x"00000000",
		2180 =>	x"00000000",
		2181 =>	x"000B0C0D",
		2182 =>	x"0E0F0000",
		2183 =>	x"10001112",
		2184 =>	x"00000000",
		2185 =>	x"00131415",
		2186 =>	x"16170800",
		2187 =>	x"00000000",
		2188 =>	x"00000000",
		2189 =>	x"00000000",
		2190 =>	x"00000000",
		2191 =>	x"00000000",
		2192 =>	x"00000000",
		2193 =>	x"00000000",
		2194 =>	x"00000000",
		2195 =>	x"00000000",
		2196 =>	x"00000000",
		2197 =>	x"00000000",
		2198 =>	x"00000000",
		2199 =>	x"00000000",
		2200 =>	x"00000000",
		2201 =>	x"00000000",
		2202 =>	x"00000000",
		2203 =>	x"00000000",
		2204 =>	x"00000000",
		2205 =>	x"00000000",
		2206 =>	x"00000000",
		2207 =>	x"00000000",
		2208 =>	x"00000000",
		2209 =>	x"00000000",
		2210 =>	x"00000000",
		2211 =>	x"00000000",
		2212 =>	x"18191A1B",
		2213 =>	x"1C1D1C1B",
		2214 =>	x"1E1F2000",
		2215 =>	x"00000000",
		2216 =>	x"30303042",
		2217 =>	x"43444515",
		2218 =>	x"2117462B",
		2219 =>	x"2C2D2E2F",
		2220 =>	x"30303030",
		2221 =>	x"30303030",
		2222 =>	x"30303030",
		2223 =>	x"30303030",
		2224 =>	x"30303030",
		2225 =>	x"30303030",
		2226 =>	x"30303030",
		2227 =>	x"30303030",
		2228 =>	x"30303030",
		2229 =>	x"30303030",
		2230 =>	x"30303030",
		2231 =>	x"30303030",
		2232 =>	x"30303030",
		2233 =>	x"30303030",
		2234 =>	x"30303030",
		2235 =>	x"30303030",
		2236 =>	x"33343536",
		2237 =>	x"37252627",
		2238 =>	x"30303030",
		2239 =>	x"30303030",
		2240 =>	x"02030405", -- IMG_16x16_rock
		2241 =>	x"06070800",
		2242 =>	x"0000090A",
		2243 =>	x"00000000",
		2244 =>	x"00000000",
		2245 =>	x"000B0C0D",
		2246 =>	x"0E0F0000",
		2247 =>	x"10001112",
		2248 =>	x"00000000",
		2249 =>	x"00131415",
		2250 =>	x"16170800",
		2251 =>	x"00000000",
		2252 =>	x"00000000",
		2253 =>	x"00000000",
		2254 =>	x"00000000",
		2255 =>	x"00000000",
		2256 =>	x"00000000",
		2257 =>	x"00000000",
		2258 =>	x"00000000",
		2259 =>	x"00000000",
		2260 =>	x"00000000",
		2261 =>	x"00000000",
		2262 =>	x"00000000",
		2263 =>	x"00000000",
		2264 =>	x"00000000",
		2265 =>	x"00000000",
		2266 =>	x"00000000",
		2267 =>	x"00000000",
		2268 =>	x"00000000",
		2269 =>	x"00000000",
		2270 =>	x"00000000",
		2271 =>	x"00000000",
		2272 =>	x"00000000",
		2273 =>	x"00000000",
		2274 =>	x"00000000",
		2275 =>	x"00000000",
		2276 =>	x"18191A1B",
		2277 =>	x"1C1D1C1B",
		2278 =>	x"1E1F2000",
		2279 =>	x"00000000",
		2280 =>	x"21174742",
		2281 =>	x"43444515",
		2282 =>	x"2117462B",
		2283 =>	x"2C2D2E2F",
		2284 =>	x"30303030",
		2285 =>	x"30303030",
		2286 =>	x"30303030",
		2287 =>	x"30313215",
		2288 =>	x"30303030",
		2289 =>	x"30303030",
		2290 =>	x"30303030",
		2291 =>	x"30303030",
		2292 =>	x"30303030",
		2293 =>	x"30303030",
		2294 =>	x"30303030",
		2295 =>	x"30303030",
		2296 =>	x"30303030",
		2297 =>	x"30303030",
		2298 =>	x"30303030",
		2299 =>	x"30303030",
		2300 =>	x"33343536",
		2301 =>	x"37252627",
		2302 =>	x"30303030",
		2303 =>	x"30303030",
		2304 =>	x"38383838", -- IMG_16x16_smoke
		2305 =>	x"38383838",
		2306 =>	x"38383838",
		2307 =>	x"38383838",
		2308 =>	x"38383800",
		2309 =>	x"00000038",
		2310 =>	x"38383838",
		2311 =>	x"38000038",
		2312 =>	x"3838003A",
		2313 =>	x"3A3A0000",
		2314 =>	x"00000038",
		2315 =>	x"003A3A00",
		2316 =>	x"38003A3A",
		2317 =>	x"3A3A003A",
		2318 =>	x"3A3A3A38",
		2319 =>	x"003A3A00",
		2320 =>	x"3800003A",
		2321 =>	x"3A3A3A3A",
		2322 =>	x"3A3A3A00",
		2323 =>	x"3A3A3A00",
		2324 =>	x"3A3A3A3A",
		2325 =>	x"3A000000",
		2326 =>	x"3A3A0000",
		2327 =>	x"3A3A0038",
		2328 =>	x"3A3A3A3A",
		2329 =>	x"003A3A3A",
		2330 =>	x"003A3A3A",
		2331 =>	x"3A3A3A00",
		2332 =>	x"383A3A00",
		2333 =>	x"3A3A3A3A",
		2334 =>	x"0000003A",
		2335 =>	x"3A3A3A00",
		2336 =>	x"3A3A3A00",
		2337 =>	x"3A3A3A3A",
		2338 =>	x"3A3A003A",
		2339 =>	x"3A3A3A00",
		2340 =>	x"003A3A3A",
		2341 =>	x"3A3A3A3A",
		2342 =>	x"3A3A003A",
		2343 =>	x"3A3A3838",
		2344 =>	x"3A3A3A3A",
		2345 =>	x"3A3A3A3A",
		2346 =>	x"3A3A003A",
		2347 =>	x"00000038",
		2348 =>	x"38003A3A",
		2349 =>	x"3A3A3A3A",
		2350 =>	x"3A3A003A",
		2351 =>	x"3A3A3A38",
		2352 =>	x"38003A3A",
		2353 =>	x"3A3A3A3A",
		2354 =>	x"003A3A3A",
		2355 =>	x"3A3A0038",
		2356 =>	x"003A3A3A",
		2357 =>	x"3A003A3A",
		2358 =>	x"003A3A3A",
		2359 =>	x"3A3A0038",
		2360 =>	x"00000000",
		2361 =>	x"00003A3A",
		2362 =>	x"003A3A3A",
		2363 =>	x"3A000038",
		2364 =>	x"38383838",
		2365 =>	x"38380000",
		2366 =>	x"38380000",
		2367 =>	x"00383838",


--			***** MAP *****


		2368 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2369 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2370 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2371 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2372 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2373 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2374 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2375 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2376 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2377 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2378 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2379 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2380 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2381 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2382 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2383 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2384 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2385 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2386 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2387 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2388 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2389 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2390 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2391 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2392 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2393 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2394 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2395 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2396 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2397 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2398 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2399 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2400 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2401 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2402 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2403 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2404 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2405 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2406 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2407 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2408 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2409 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2410 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2411 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2412 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2413 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2414 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2415 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2416 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2417 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2418 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2419 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2420 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2421 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2422 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2423 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2424 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2425 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2426 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2427 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2428 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2429 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2430 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2431 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2432 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2433 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2434 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2435 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2436 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2437 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2438 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2439 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2440 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2441 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2442 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2443 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2444 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2445 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2446 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2447 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2448 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2449 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2450 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2451 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2452 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2453 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2454 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2455 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2456 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2457 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2458 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2459 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2460 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2461 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2462 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2463 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2464 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2465 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2466 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2467 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2468 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2469 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2470 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2471 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2472 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2473 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2474 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2475 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2476 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2477 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2478 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2479 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2480 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2481 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2482 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2483 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2484 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2485 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2486 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2487 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2488 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2489 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2490 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2491 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2492 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2493 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2494 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2495 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2496 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2497 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2498 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2499 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2500 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2501 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2502 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2503 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2504 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2505 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2506 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2507 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2508 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2509 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2510 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2511 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2512 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2513 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2514 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2515 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2516 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2517 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2518 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2519 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2520 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2521 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2522 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2523 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2524 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2525 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2526 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2527 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2528 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2529 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2530 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2531 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2532 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2533 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2534 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2535 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2536 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2537 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2538 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2539 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2540 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2541 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2542 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2543 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2544 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2545 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2546 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2547 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2548 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2549 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2550 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2551 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2552 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2553 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2554 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2555 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2556 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2557 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2558 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2559 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2560 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2561 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2562 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2563 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2564 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2565 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2566 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2567 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2568 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2569 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2570 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2571 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2572 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2573 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2574 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2575 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2576 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2577 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2578 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2579 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2580 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2581 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2582 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2583 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2584 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2585 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2586 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2587 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2588 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2589 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2590 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2591 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2592 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2593 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2594 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2595 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2596 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2597 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2598 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2599 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2600 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2601 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2602 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2603 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2604 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2605 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2606 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2607 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2608 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2609 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2610 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2611 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2612 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2613 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2614 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2615 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2616 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2617 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2618 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2619 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2620 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2621 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2622 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2623 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2624 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2625 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2626 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2627 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2628 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2629 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2630 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2631 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2632 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2633 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2634 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2635 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2636 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2637 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2638 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2639 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2640 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2641 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2642 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2643 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2644 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2645 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2646 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2647 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2648 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2649 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2650 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2651 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2652 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2653 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2654 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2655 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2656 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2657 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2658 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2659 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2660 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2661 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2662 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2663 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2664 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2665 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2666 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2667 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2668 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2669 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2670 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2671 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2672 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2673 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2674 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2675 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2676 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2677 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2678 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2679 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2680 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2681 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2682 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2683 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2684 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2685 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2686 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2687 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2688 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2689 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2690 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2691 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2692 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2693 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2694 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2695 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2696 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2697 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2698 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2699 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2700 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2701 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2702 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2703 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2704 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2705 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2706 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2707 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2708 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2709 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2710 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2711 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2712 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2713 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2714 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2715 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2716 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2717 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2718 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2719 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2720 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2721 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2722 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2723 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2724 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2725 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2726 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2727 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2728 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2729 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2730 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2731 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2732 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2733 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2734 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2735 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2736 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2737 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2738 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2739 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2740 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2741 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2742 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2743 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2744 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2745 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2746 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2747 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2748 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2749 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2750 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2751 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2752 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2753 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2754 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2755 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2756 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2757 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2758 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2759 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2760 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2761 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2762 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2763 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2764 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2765 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2766 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2767 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2768 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2769 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2770 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2771 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2772 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2773 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2774 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2775 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2776 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2777 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2778 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2779 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2780 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2781 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2782 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2783 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2784 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2785 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2786 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2787 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2788 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2789 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2790 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2791 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2792 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2793 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2794 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2795 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2796 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2797 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2798 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2799 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2800 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2801 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2802 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2803 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2804 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2805 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2806 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2807 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2808 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2809 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2810 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2811 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2812 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2813 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2814 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2815 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2816 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2817 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2818 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2819 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2820 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2821 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2822 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2823 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2824 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2825 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2826 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2827 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2828 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2829 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2830 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2831 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2832 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2833 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2834 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2835 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2836 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2837 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2838 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2839 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2840 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2841 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2842 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2843 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2844 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2845 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2846 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2847 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2848 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2849 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2850 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2851 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2852 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2853 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2854 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2855 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2856 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2857 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2858 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2859 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2860 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2861 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2862 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2863 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2864 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2865 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2866 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2867 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2868 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2869 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2870 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2871 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2872 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2873 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2874 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2875 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2876 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2877 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2878 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2879 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2880 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2881 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2882 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2883 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2884 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2885 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2886 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2887 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2888 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2889 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2890 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2891 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2892 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2893 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2894 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2895 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2896 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2897 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2898 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2899 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2900 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2901 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2902 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2903 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2904 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2905 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2906 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2907 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2908 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2909 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2910 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2911 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2912 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2913 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2914 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2915 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2916 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2917 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2918 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2919 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2920 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2921 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2922 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2923 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2924 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2925 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2926 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2927 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2928 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2929 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2930 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2931 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2932 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2933 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2934 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2935 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2936 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2937 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2938 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2939 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2940 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2941 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2942 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2943 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2944 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2945 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2946 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2947 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2948 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2949 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2950 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2951 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2952 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2953 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2954 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2955 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2956 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2957 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2958 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2959 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2960 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2961 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2962 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2963 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2964 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2965 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2966 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2967 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2968 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2969 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2970 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2971 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2972 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2973 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2974 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2975 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2976 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2977 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2978 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2979 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2980 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2981 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2982 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2983 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2984 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2985 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2986 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2987 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2988 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2989 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2990 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2991 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2992 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2993 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2994 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2995 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2996 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2997 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2998 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2999 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3000 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3001 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3002 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3003 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3004 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3005 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3006 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3007 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3008 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3009 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3010 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3011 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3012 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3013 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3014 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3015 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3016 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3017 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3018 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3019 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3020 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3021 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3022 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3023 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3024 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3025 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3026 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3027 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3028 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3029 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3030 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3031 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3032 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3033 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3034 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3035 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3036 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3037 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3038 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3039 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3040 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3041 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3042 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3043 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3044 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3045 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3046 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3047 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3048 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3049 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3050 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3051 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3052 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3053 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3054 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3055 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3056 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3057 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3058 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3059 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3060 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3061 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3062 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3063 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3064 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3065 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3066 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3067 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3068 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3069 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3070 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3071 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3072 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3073 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3074 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3075 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3076 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3077 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3078 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3079 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3080 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3081 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3082 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3083 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3084 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3085 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3086 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3087 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3088 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3089 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3090 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3091 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3092 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3093 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3094 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3095 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3096 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3097 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3098 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3099 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3100 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3101 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3102 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3103 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3104 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3105 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3106 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3107 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3108 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3109 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3110 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3111 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3112 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3113 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3114 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3115 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3116 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3117 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3118 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3119 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3120 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3121 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3122 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3123 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3124 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3125 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3126 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3127 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3128 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3129 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3130 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3131 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3132 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3133 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3134 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3135 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3136 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3137 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3138 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3139 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3140 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3141 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3142 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3143 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3144 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3145 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3146 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3147 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3148 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3149 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3150 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3151 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3152 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3153 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3154 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3155 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3156 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3157 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3158 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3159 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3160 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3161 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3162 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3163 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3164 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3165 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3166 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3167 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3168 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3169 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3170 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3171 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3172 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3173 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3174 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3175 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3176 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3177 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3178 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3179 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3180 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3181 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3182 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3183 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3184 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3185 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3186 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3187 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3188 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3189 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3190 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3191 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3192 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3193 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3194 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3195 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3196 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3197 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3198 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3199 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3200 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3201 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3202 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3203 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3204 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3205 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3206 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3207 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3208 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3209 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3210 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3211 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3212 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3213 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3214 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3215 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3216 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3217 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3218 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3219 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3220 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3221 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3222 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3223 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3224 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3225 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3226 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3227 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3228 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3229 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3230 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3231 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3232 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3233 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3234 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3235 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3236 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3237 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3238 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3239 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3240 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3241 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3242 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3243 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3244 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3245 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3246 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3247 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3248 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3249 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3250 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3251 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3252 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3253 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3254 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3255 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3256 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3257 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3258 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3259 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3260 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3261 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3262 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3263 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3264 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3265 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3266 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3267 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3268 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3269 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3270 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3271 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3272 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3273 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3274 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3275 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3276 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3277 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3278 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3279 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3280 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3281 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3282 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3283 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3284 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3285 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3286 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3287 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3288 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3289 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3290 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3291 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3292 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3293 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3294 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3295 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3296 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3297 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3298 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3299 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3300 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3301 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3302 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3303 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3304 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3305 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3306 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3307 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3308 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3309 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3310 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3311 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3312 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3313 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3314 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3315 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3316 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3317 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3318 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3319 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3320 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3321 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3322 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3323 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3324 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3325 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3326 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3327 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3328 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3329 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3330 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3331 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3332 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3333 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3334 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3335 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3336 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3337 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3338 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3339 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3340 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3341 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3342 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3343 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3344 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3345 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3346 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3347 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3348 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3349 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3350 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3351 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3352 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3353 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3354 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3355 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3356 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3357 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3358 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3359 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3360 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3361 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3362 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3363 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3364 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3365 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3366 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3367 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3368 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3369 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3370 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3371 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3372 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3373 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3374 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3375 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3376 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3377 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3378 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3379 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3380 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3381 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3382 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3383 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3384 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3385 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3386 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3387 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3388 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3389 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3390 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3391 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3392 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3393 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3394 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3395 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3396 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3397 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3398 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3399 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3400 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3401 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3402 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3403 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3404 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3405 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3406 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3407 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3408 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3409 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3410 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3411 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3412 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3413 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3414 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3415 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3416 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3417 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3418 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3419 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3420 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3421 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3422 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3423 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3424 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3425 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3426 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3427 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3428 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3429 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3430 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3431 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3432 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3433 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3434 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3435 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3436 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3437 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3438 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3439 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3440 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3441 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3442 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3443 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3444 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3445 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3446 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3447 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3448 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3449 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3450 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3451 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3452 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3453 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3454 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3455 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3456 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3457 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3458 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3459 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3460 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3461 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3462 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3463 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3464 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3465 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3466 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3467 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3468 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3469 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3470 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3471 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3472 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3473 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3474 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3475 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3476 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3477 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3478 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3479 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3480 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3481 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3482 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3483 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3484 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3485 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3486 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3487 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3488 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3489 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3490 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3491 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3492 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3493 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3494 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3495 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3496 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3497 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3498 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3499 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3500 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3501 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3502 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3503 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3504 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3505 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3506 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3507 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3508 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3509 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3510 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3511 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3512 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3513 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3514 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3515 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3516 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3517 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3518 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3519 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3520 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3521 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3522 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3523 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3524 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3525 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3526 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3527 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3528 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3529 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3530 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3531 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3532 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3533 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3534 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3535 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3536 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3537 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3538 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3539 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3540 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3541 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3542 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3543 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3544 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3545 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3546 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3547 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3548 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3549 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3550 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3551 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3552 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3553 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3554 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3555 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3556 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3557 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3558 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3559 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3560 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3561 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3562 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3563 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3564 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3565 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3566 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3567 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3568 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3569 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3570 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3571 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3572 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3573 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3574 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3575 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3576 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3577 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3578 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3579 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3580 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3581 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3582 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3583 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3584 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3585 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3586 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3587 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3588 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3589 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3590 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3591 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3592 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3593 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3594 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3595 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3596 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3597 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3598 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3599 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3600 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3601 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3602 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3603 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3604 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3605 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3606 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3607 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3608 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3609 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3610 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3611 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3612 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3613 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3614 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3615 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3616 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3617 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3618 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3619 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3620 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3621 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3622 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3623 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3624 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3625 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3626 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3627 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3628 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3629 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3630 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3631 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3632 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3633 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3634 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3635 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3636 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3637 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3638 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;