
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER
-- DATE: Thu May 24 09:52:20 2018

	signal mem : ram_t := (
	

--			***** COLOR PALLETE *****


		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00277FFF", -- R: 255 G: 127 B: 39
		2 =>	x"00433A5C", -- R: 92 G: 58 B: 67
		3 =>	x"0050726F", -- R: 111 G: 114 B: 80
		4 =>	x"00677261", -- R: 97 G: 114 B: 103
		5 =>	x"006D4461", -- R: 97 G: 68 B: 109
		6 =>	x"00746100", -- R: 0 G: 97 B: 116
		7 =>	x"00FDFDFD", -- R: 253 G: 253 B: 253
		8 =>	x"00FD0000", -- R: 0 G: 0 B: 253
		9 =>	x"003A04D7", -- R: 215 G: 4 B: 58
		10 =>	x"0013549B", -- R: 155 G: 84 B: 19
		11 =>	x"00000C98", -- R: 152 G: 12 B: 0
		12 =>	x"009B5B00", -- R: 0 G: 91 B: 155
		13 =>	x"0060A05B", -- R: 91 G: 160 B: 96
		14 =>	x"0000F424", -- R: 36 G: 244 B: 0
		15 =>	x"00850F40", -- R: 64 G: 15 B: 133
		16 =>	x"0028AF5B", -- R: 91 G: 175 B: 40
		17 =>	x"00006872", -- R: 114 G: 104 B: 0
		18 =>	x"005B0078", -- R: 120 G: 0 B: 91
		19 =>	x"0057870F", -- R: 15 G: 135 B: 87
		20 =>	x"00810000", -- R: 0 G: 0 B: 129
		21 =>	x"00000200", -- R: 0 G: 2 B: 0
		22 =>	x"0000001F", -- R: 31 G: 0 B: 0
		23 =>	x"000D0000", -- R: 0 G: 0 B: 13
		24 =>	x"0000FDFD", -- R: 253 G: 253 B: 0
		25 =>	x"00FDFD41", -- R: 65 G: 253 B: 253
		26 =>	x"004C4C55", -- R: 85 G: 76 B: 76
		27 =>	x"00534552", -- R: 82 G: 69 B: 83
		28 =>	x"00535052", -- R: 82 G: 80 B: 83
		29 =>	x"004F4649", -- R: 73 G: 70 B: 79
		30 =>	x"004C453D", -- R: 61 G: 69 B: 76
		31 =>	x"00020000", -- R: 0 G: 0 B: 2
		32 =>	x"00000F00", -- R: 0 G: 15 B: 0
		33 =>	x"0000000C", -- R: 12 G: 0 B: 0
		34 =>	x"00FD4144", -- R: 68 G: 65 B: 253
		35 =>	x"00564958", -- R: 88 G: 73 B: 86
		36 =>	x"00455F4C", -- R: 76 G: 95 B: 69
		37 =>	x"00414E47", -- R: 71 G: 78 B: 65
		38 =>	x"003D656E", -- R: 110 G: 101 B: 61
		39 =>	x"00FDFD00", -- R: 0 G: 253 B: 253
		40 =>	x"00003606", -- R: 6 G: 54 B: 0
		41 =>	x"00D71D56", -- R: 86 G: 29 B: 215
		42 =>	x"009B000D", -- R: 13 G: 0 B: 155
		43 =>	x"006F6F6C", -- R: 108 G: 111 B: 111
		44 =>	x"00735C41", -- R: 65 G: 92 B: 115
		45 =>	x"00647669", -- R: 105 G: 118 B: 100
		46 =>	x"00736F72", -- R: 114 G: 111 B: 115
		47 =>	x"00203230", -- R: 48 G: 50 B: 32
		48 =>	x"0031375C", -- R: 92 G: 55 B: 49
		49 =>	x"003406D7", -- R: 215 G: 6 B: 52
		50 =>	x"001F509B", -- R: 155 G: 80 B: 31
		51 =>	x"00000DB8", -- R: 184 G: 13 B: 0
		52 =>	x"00AE5B00", -- R: 0 G: 91 B: 174
		53 =>	x"0068AF5B", -- R: 91 G: 175 B: 104
		54 =>	x"00007857", -- R: 87 G: 120 B: 0
		55 =>	x"00870F81", -- R: 129 G: 15 B: 135
		56 =>	x"00414456", -- R: 86 G: 68 B: 65
		57 =>	x"0049534F", -- R: 79 G: 83 B: 73
		58 =>	x"00525F32", -- R: 50 G: 95 B: 82
		59 =>	x"00303137", -- R: 55 G: 49 B: 48
		60 =>	x"005F4449", -- R: 73 G: 68 B: 95
		61 =>	x"00523D43", -- R: 67 G: 61 B: 82
		62 =>	x"003A5C50", -- R: 80 G: 92 B: 58
		63 =>	x"00726F67", -- R: 103 G: 111 B: 114
		64 =>	x"0072616D", -- R: 109 G: 97 B: 114
		65 =>	x"00204669", -- R: 105 G: 70 B: 32
		66 =>	x"006C6573", -- R: 115 G: 101 B: 108
		67 =>	x"00202878", -- R: 120 G: 40 B: 32
		68 =>	x"00383629", -- R: 41 G: 54 B: 56
		69 =>	x"005C496E", -- R: 110 G: 73 B: 92
		70 =>	x"0074656C", -- R: 108 G: 101 B: 116
		71 =>	x"00535754", -- R: 84 G: 87 B: 83
		72 =>	x"00DDDDDD", -- R: 221 G: 221 B: 221
		73 =>	x"00000032", -- R: 50 G: 0 B: 0
		74 =>	x"0006D719", -- R: 25 G: 215 B: 6
		75 =>	x"005D9B00", -- R: 0 G: 155 B: 93
		76 =>	x"00091871", -- R: 113 G: 24 B: 9
		77 =>	x"005B0028", -- R: 40 G: 0 B: 91
		78 =>	x"00AF5B00", -- R: 0 G: 91 B: 175
		79 =>	x"00785787", -- R: 135 G: 87 B: 120
		80 =>	x"000F8100", -- R: 0 G: 129 B: 15
		81 =>	x"00000002", -- R: 2 G: 0 B: 0
		82 =>	x"00430000", -- R: 0 G: 0 B: 67
		83 =>	x"00000B00", -- R: 0 G: 11 B: 0
		84 =>	x"000000FD", -- R: 253 G: 0 B: 0
		85 =>	x"0069006E", -- R: 110 G: 0 B: 105
		86 =>	x"00006400", -- R: 0 G: 100 B: 0
		87 =>	x"006F0077", -- R: 119 G: 0 B: 111
		88 =>	x"00007300", -- R: 0 G: 115 B: 0
		89 =>	x"005C0072", -- R: 114 G: 0 B: 92
		90 =>	x"00006500", -- R: 0 G: 101 B: 0
		91 =>	x"00730063", -- R: 99 G: 0 B: 115
		92 =>	x"00006100", -- R: 0 G: 97 B: 0
		93 =>	x"00630068", -- R: 104 G: 0 B: 99
		94 =>	x"0000003F", -- R: 63 G: 0 B: 0
		95 =>	x"0006D615", -- R: 21 G: 214 B: 6
		96 =>	x"00589B00", -- R: 0 G: 155 B: 88
		97 =>	x"0000D8AC", -- R: 172 G: 216 B: 0
		98 =>	x"005B00C4", -- R: 196 G: 0 B: 91
		99 =>	x"00005700", -- R: 0 G: 87 B: 0
		100 =>	x"003806D7", -- R: 215 G: 6 B: 56
		101 =>	x"0013589B", -- R: 155 G: 88 B: 19
		102 =>	x"00000C03", -- R: 3 G: 12 B: 0
		103 =>	x"00001000", -- R: 0 G: 16 B: 0
		104 =>	x"00280010", -- R: 16 G: 0 B: 40
		105 =>	x"0000DDDD", -- R: 221 G: 221 B: 0
		106 =>	x"00DDDD3A", -- R: 58 G: 221 B: 221
		107 =>	x"0006D711", -- R: 17 G: 215 B: 6
		108 =>	x"005A9B00", -- R: 0 G: 155 B: 90
		109 =>	x"00084300", -- R: 0 G: 67 B: 8
		110 =>	x"003A005C", -- R: 92 G: 0 B: 58
		111 =>	x"003A06D7", -- R: 215 G: 6 B: 58
		112 =>	x"0011459B", -- R: 155 G: 69 B: 17
		113 =>	x"00000C01", -- R: 1 G: 12 B: 0
		114 =>	x"0000FFFF", -- R: 255 G: 255 B: 0
		115 =>	x"00FFFF00", -- R: 0 G: 255 B: 255
		116 =>	x"0068000F", -- R: 15 G: 0 B: 104
		117 =>	x"0000C800", -- R: 0 G: 200 B: 0
		118 =>	x"000F00F0", -- R: 240 G: 0 B: 15
		119 =>	x"000050AE", -- R: 174 G: 80 B: 0
		120 =>	x"005B00DD", -- R: 221 G: 0 B: 91
		121 =>	x"00000009", -- R: 9 G: 0 B: 0
		122 =>	x"0080AD5B", -- R: 91 G: 173 B: 128
		123 =>	x"00000001", -- R: 1 G: 0 B: 0
		124 =>	x"00004000", -- R: 0 G: 64 B: 0
		125 =>	x"00000035", -- R: 53 G: 0 B: 0
		126 =>	x"00003200", -- R: 0 G: 50 B: 0
		127 =>	x"00430036", -- R: 54 G: 0 B: 67
		128 =>	x"00003400", -- R: 0 G: 52 B: 0
		129 =>	x"00420037", -- R: 55 G: 0 B: 66
		130 =>	x"00004500", -- R: 0 G: 69 B: 0
		131 =>	x"00000100", -- R: 0 G: 1 B: 0
		132 =>	x"002706D7", -- R: 215 G: 6 B: 39
		133 =>	x"000C579B", -- R: 155 G: 87 B: 12
		134 =>	x"00000ACE", -- R: 206 G: 10 B: 0
		135 =>	x"00020019", -- R: 25 G: 0 B: 2
		136 =>	x"00000040", -- R: 64 G: 0 B: 0
		137 =>	x"00AA5B00", -- R: 0 G: 91 B: 170
		138 =>	x"003506D7", -- R: 215 G: 6 B: 53
		139 =>	x"001E5B9B", -- R: 155 G: 91 B: 30
		140 =>	x"00000A3E", -- R: 62 G: 10 B: 0
		141 =>	x"00010001", -- R: 1 G: 0 B: 1
		142 =>	x"0038AD5B", -- R: 91 G: 173 B: 56
		143 =>	x"00005000", -- R: 0 G: 80 B: 0
		144 =>	x"00000039", -- R: 57 G: 0 B: 0
		145 =>	x"0006D613", -- R: 19 G: 214 B: 6
		146 =>	x"000020A7", -- R: 167 G: 32 B: 0
		147 =>	x"005B00A0", -- R: 160 G: 0 B: 91
		148 =>	x"007F7F7F", -- R: 127 G: 127 B: 127
		149 =>	x"00FF0000", -- R: 0 G: 0 B: 255
		150 =>	x"004798FF", -- R: 255 G: 152 B: 71
		151 =>	x"000000FF", -- R: 255 G: 0 B: 0
		152 =>	x"00007F00", -- R: 0 G: 127 B: 0
		153 =>	x"004C4C4C", -- R: 76 G: 76 B: 76
		154 =>	x"007F007F", -- R: 127 G: 0 B: 127
		155 =>	x"0000007F", -- R: 127 G: 0 B: 0
		156 =>	x"00007F82", -- R: 130 G: 127 B: 0
		157 =>	x"00666666", -- R: 102 G: 102 B: 102
		158 =>	x"009800FF", -- R: 255 G: 0 B: 152
		159 =>	x"009800A4", -- R: 164 G: 0 B: 152
		160 =>	x"00980000", -- R: 0 G: 0 B: 152
		161 =>	x"005480D7", -- R: 215 G: 128 B: 84
		162 =>	x"00862138", -- R: 56 G: 33 B: 134
		163 =>	x"00990000", -- R: 0 G: 0 B: 153
		164 =>	x"00862136", -- R: 54 G: 33 B: 134
		165 =>	x"00980124", -- R: 36 G: 1 B: 152
		166 =>	x"00980095", -- R: 149 G: 0 B: 152
		167 =>	x"009800A5", -- R: 165 G: 0 B: 152
		168 =>	x"00980094", -- R: 148 G: 0 B: 152
		169 =>	x"009800DF", -- R: 223 G: 0 B: 152
		170 =>	x"009800A7", -- R: 167 G: 0 B: 152
		171 =>	x"0098016B", -- R: 107 G: 1 B: 152
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
		255 =>	x"00000000", -- Unused


--			***** 16x16 IMAGES *****


		256 =>	x"01010101", -- IMG_16x16_background
		257 =>	x"01010101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01010101",
		261 =>	x"01010101",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01010101",
		265 =>	x"01010101",
		266 =>	x"01010101",
		267 =>	x"01010101",
		268 =>	x"01010101",
		269 =>	x"01010101",
		270 =>	x"01010101",
		271 =>	x"01010101",
		272 =>	x"01010101",
		273 =>	x"01010101",
		274 =>	x"01010101",
		275 =>	x"01010101",
		276 =>	x"01010101",
		277 =>	x"01010101",
		278 =>	x"01010101",
		279 =>	x"01010101",
		280 =>	x"01010101",
		281 =>	x"01010101",
		282 =>	x"01010101",
		283 =>	x"01010101",
		284 =>	x"01010101",
		285 =>	x"01010101",
		286 =>	x"01010101",
		287 =>	x"01010101",
		288 =>	x"01010101",
		289 =>	x"01010101",
		290 =>	x"01010101",
		291 =>	x"01010101",
		292 =>	x"01010101",
		293 =>	x"01010101",
		294 =>	x"01010101",
		295 =>	x"01010101",
		296 =>	x"01010101",
		297 =>	x"01010101",
		298 =>	x"01010101",
		299 =>	x"01010101",
		300 =>	x"01010101",
		301 =>	x"01010101",
		302 =>	x"01010101",
		303 =>	x"01010101",
		304 =>	x"01010101",
		305 =>	x"01010101",
		306 =>	x"01010101",
		307 =>	x"01010101",
		308 =>	x"01010101",
		309 =>	x"01010101",
		310 =>	x"01010101",
		311 =>	x"01010101",
		312 =>	x"01010101",
		313 =>	x"01010101",
		314 =>	x"01010101",
		315 =>	x"01010101",
		316 =>	x"01010101",
		317 =>	x"01010101",
		318 =>	x"01010101",
		319 =>	x"01010101",
		320 =>	x"02030405", -- IMG_16x16_bang
		321 =>	x"06070800",
		322 =>	x"090A0B0C",
		323 =>	x"0D0E0F00",
		324 =>	x"10111213",
		325 =>	x"14151600",
		326 =>	x"1718191A",
		327 =>	x"1B1C1D1E",
		328 =>	x"1F202100",
		329 =>	x"07222324",
		330 =>	x"25261827",
		331 =>	x"0028292A",
		332 =>	x"2B2C2D2E",
		333 =>	x"2F301827",
		334 =>	x"31323334",
		335 =>	x"35363700",
		336 =>	x"38393A3B",
		337 =>	x"3C3D3E3F",
		338 =>	x"40414243",
		339 =>	x"44454647",
		340 =>	x"4800494A",
		341 =>	x"4B4C4D4E",
		342 =>	x"4F505100",
		343 =>	x"52535407",
		344 =>	x"55565758",
		345 =>	x"595A5B5C",
		346 =>	x"5D5A5E5F",
		347 =>	x"60616263",
		348 =>	x"64656600",
		349 =>	x"00000067",
		350 =>	x"68696A6B",
		351 =>	x"6C6D6E63",
		352 =>	x"6F707100",
		353 =>	x"00727320",
		354 =>	x"74757620",
		355 =>	x"00777848",
		356 =>	x"00000000",
		357 =>	x"00000000",
		358 =>	x"00000000",
		359 =>	x"00000069",
		360 =>	x"00000000",
		361 =>	x"00000000",
		362 =>	x"00000000",
		363 =>	x"00000000",
		364 =>	x"79000000",
		365 =>	x"00000000",
		366 =>	x"00000000",
		367 =>	x"00000000",
		368 =>	x"7A007B00",
		369 =>	x"007C7D7E",
		370 =>	x"7F808182",
		371 =>	x"00150083",
		372 =>	x"00000000",
		373 =>	x"00150069",
		374 =>	x"84858600",
		375 =>	x"87008889",
		376 =>	x"8A8B8C00",
		377 =>	x"8D838889",
		378 =>	x"8E000000",
		379 =>	x"008F0000",
		380 =>	x"07089091",
		381 =>	x"60929334",
		382 =>	x"00000000",
		383 =>	x"00004848",
		384 =>	x"00000000", -- IMG_16x16_car_blue
		385 =>	x"00000000",
		386 =>	x"00000000",
		387 =>	x"00000000",
		388 =>	x"00009494",
		389 =>	x"94000000",
		390 =>	x"00000000",
		391 =>	x"00000000",
		392 =>	x"00009494",
		393 =>	x"94000095",
		394 =>	x"00000000",
		395 =>	x"00000000",
		396 =>	x"00000094",
		397 =>	x"00000095",
		398 =>	x"95000000",
		399 =>	x"00000000",
		400 =>	x"00009595",
		401 =>	x"95959595",
		402 =>	x"95950000",
		403 =>	x"94949400",
		404 =>	x"00949495",
		405 =>	x"95959595",
		406 =>	x"95959595",
		407 =>	x"94949400",
		408 =>	x"00949494",
		409 =>	x"94727272",
		410 =>	x"95959595",
		411 =>	x"00940000",
		412 =>	x"00009595",
		413 =>	x"95727272",
		414 =>	x"72959595",
		415 =>	x"95959500",
		416 =>	x"00009595",
		417 =>	x"95727272",
		418 =>	x"72959595",
		419 =>	x"95959500",
		420 =>	x"00949494",
		421 =>	x"94727272",
		422 =>	x"95959595",
		423 =>	x"00940000",
		424 =>	x"00949495",
		425 =>	x"95959595",
		426 =>	x"95959595",
		427 =>	x"94949400",
		428 =>	x"00009595",
		429 =>	x"95959595",
		430 =>	x"95950000",
		431 =>	x"94949400",
		432 =>	x"00000094",
		433 =>	x"00000095",
		434 =>	x"95000000",
		435 =>	x"00000000",
		436 =>	x"00009494",
		437 =>	x"94000095",
		438 =>	x"00000000",
		439 =>	x"00000000",
		440 =>	x"00009494",
		441 =>	x"94000000",
		442 =>	x"00000000",
		443 =>	x"00000000",
		444 =>	x"00000000",
		445 =>	x"00000000",
		446 =>	x"00000000",
		447 =>	x"00000000",
		448 =>	x"96969696", -- IMG_16x16_car_red
		449 =>	x"96969696",
		450 =>	x"96969696",
		451 =>	x"96969696",
		452 =>	x"96960000",
		453 =>	x"00969696",
		454 =>	x"96969696",
		455 =>	x"96969696",
		456 =>	x"96960000",
		457 =>	x"00969697",
		458 =>	x"96969696",
		459 =>	x"96969696",
		460 =>	x"96969600",
		461 =>	x"96969697",
		462 =>	x"97969696",
		463 =>	x"96969696",
		464 =>	x"96969797",
		465 =>	x"97979797",
		466 =>	x"97979696",
		467 =>	x"00000096",
		468 =>	x"96000097",
		469 =>	x"97979797",
		470 =>	x"97979797",
		471 =>	x"00000096",
		472 =>	x"96000000",
		473 =>	x"00727272",
		474 =>	x"97979797",
		475 =>	x"96009696",
		476 =>	x"96969797",
		477 =>	x"97727272",
		478 =>	x"72979797",
		479 =>	x"97979796",
		480 =>	x"96969797",
		481 =>	x"97727272",
		482 =>	x"72979797",
		483 =>	x"97979796",
		484 =>	x"96000000",
		485 =>	x"00727272",
		486 =>	x"97979797",
		487 =>	x"96009696",
		488 =>	x"96000097",
		489 =>	x"97979797",
		490 =>	x"97979797",
		491 =>	x"00000096",
		492 =>	x"96969797",
		493 =>	x"97979797",
		494 =>	x"97979696",
		495 =>	x"00000096",
		496 =>	x"96969600",
		497 =>	x"96969697",
		498 =>	x"97969696",
		499 =>	x"96969696",
		500 =>	x"96960000",
		501 =>	x"00969697",
		502 =>	x"96969696",
		503 =>	x"96969696",
		504 =>	x"96960000",
		505 =>	x"00969696",
		506 =>	x"96969696",
		507 =>	x"96969696",
		508 =>	x"96969696",
		509 =>	x"96969696",
		510 =>	x"96969696",
		511 =>	x"96969696",
		512 =>	x"01010101", -- IMG_16x16_flag
		513 =>	x"01010101",
		514 =>	x"01010101",
		515 =>	x"01010101",
		516 =>	x"01017272",
		517 =>	x"01010101",
		518 =>	x"01010101",
		519 =>	x"01010101",
		520 =>	x"01017272",
		521 =>	x"72720101",
		522 =>	x"01010101",
		523 =>	x"01010101",
		524 =>	x"01017272",
		525 =>	x"72727272",
		526 =>	x"01010101",
		527 =>	x"01010101",
		528 =>	x"01017272",
		529 =>	x"72727272",
		530 =>	x"72720101",
		531 =>	x"01010101",
		532 =>	x"01017272",
		533 =>	x"72727272",
		534 =>	x"72727272",
		535 =>	x"01010101",
		536 =>	x"01017272",
		537 =>	x"72727272",
		538 =>	x"72720101",
		539 =>	x"01010101",
		540 =>	x"01017272",
		541 =>	x"72727272",
		542 =>	x"01010101",
		543 =>	x"01010101",
		544 =>	x"01017272",
		545 =>	x"72720101",
		546 =>	x"01010101",
		547 =>	x"01010101",
		548 =>	x"01017272",
		549 =>	x"01010101",
		550 =>	x"01010101",
		551 =>	x"01010101",
		552 =>	x"01017272",
		553 =>	x"01010101",
		554 =>	x"01010101",
		555 =>	x"01010101",
		556 =>	x"01017272",
		557 =>	x"01010101",
		558 =>	x"01010101",
		559 =>	x"01010101",
		560 =>	x"01017272",
		561 =>	x"01010101",
		562 =>	x"01010101",
		563 =>	x"01010101",
		564 =>	x"01727272",
		565 =>	x"72010101",
		566 =>	x"01010101",
		567 =>	x"01010101",
		568 =>	x"01727272",
		569 =>	x"72010101",
		570 =>	x"01010101",
		571 =>	x"01010101",
		572 =>	x"01010101",
		573 =>	x"01010101",
		574 =>	x"01010101",
		575 =>	x"01010101",
		576 =>	x"98989898", -- IMG_16x16_map_element_00
		577 =>	x"98989998",
		578 =>	x"99999898",
		579 =>	x"98989898",
		580 =>	x"98989898",
		581 =>	x"9A9B9B9A",
		582 =>	x"9B9A9B99",
		583 =>	x"98989898",
		584 =>	x"9898999B",
		585 =>	x"9A9B9B9A",
		586 =>	x"9C9D9B9B",
		587 =>	x"98989898",
		588 =>	x"98989A9B",
		589 =>	x"9B9B9A9A",
		590 =>	x"9B9B9A9A",
		591 =>	x"9B9B9898",
		592 =>	x"98999B9B",
		593 =>	x"9B9B9A9A",
		594 =>	x"9B979A9A",
		595 =>	x"9A999998",
		596 =>	x"999A9A9B",
		597 =>	x"9B979A9A",
		598 =>	x"9B979A9B",
		599 =>	x"9B9B9B99",
		600 =>	x"999B9B9B",
		601 =>	x"9B9B9B9A",
		602 =>	x"9B9B9B97",
		603 =>	x"979B9B99",
		604 =>	x"999C9A9A",
		605 =>	x"9B9A9A99",
		606 =>	x"9A9A9B9A",
		607 =>	x"979B9999",
		608 =>	x"999B9B9C",
		609 =>	x"9B9B9B9B",
		610 =>	x"9B9B9B97",
		611 =>	x"9B9B9B99",
		612 =>	x"999B9B9B",
		613 =>	x"9B9C9B9A",
		614 =>	x"9B9B9A9B",
		615 =>	x"9A9B9A99",
		616 =>	x"999A9B9B",
		617 =>	x"9B9B9A9B",
		618 =>	x"979A9B9B",
		619 =>	x"9A999A99",
		620 =>	x"989B9B9A",
		621 =>	x"9A9A9A9B",
		622 =>	x"9B9A9A9B",
		623 =>	x"9A9A9998",
		624 =>	x"98989A9B",
		625 =>	x"9B9A9B9B",
		626 =>	x"9A9A9A9B",
		627 =>	x"9B9B9998",
		628 =>	x"9898999C",
		629 =>	x"9B9A9C9B",
		630 =>	x"9A9A9B9B",
		631 =>	x"9A999898",
		632 =>	x"98989898",
		633 =>	x"999B9C9C",
		634 =>	x"9B979998",
		635 =>	x"98989898",
		636 =>	x"98989898",
		637 =>	x"98989999",
		638 =>	x"99999898",
		639 =>	x"98989898",
		640 =>	x"9E9E9E9E", -- IMG_16x16_map_element_01
		641 =>	x"9E9E9E9E",
		642 =>	x"9E9E9E9E",
		643 =>	x"9E9E9FA0",
		644 =>	x"9E9E9E9E",
		645 =>	x"9E9E9E9E",
		646 =>	x"9E9E9E9E",
		647 =>	x"9E9E9FA0",
		648 =>	x"9E9E9E9E",
		649 =>	x"9E9E9E9E",
		650 =>	x"9E9E9E9E",
		651 =>	x"9E9E9FA0",
		652 =>	x"9E9E9E9E",
		653 =>	x"9E9E9E9E",
		654 =>	x"9E9E9E9E",
		655 =>	x"9E9E9FA0",
		656 =>	x"9E9E9E9E",
		657 =>	x"9E9E9E9E",
		658 =>	x"9E9E9E9E",
		659 =>	x"9E9E9FA0",
		660 =>	x"9E9E9E9E",
		661 =>	x"9E9E9E9E",
		662 =>	x"9E9E9E9E",
		663 =>	x"9E9E9FA0",
		664 =>	x"9E9E9E9E",
		665 =>	x"9E9E9E9E",
		666 =>	x"9E9E9E9E",
		667 =>	x"9E9E9FA0",
		668 =>	x"9E9E9E9E",
		669 =>	x"9E9E9E9E",
		670 =>	x"9E9E9E9E",
		671 =>	x"9E9E9FA0",
		672 =>	x"9E9E9E9E",
		673 =>	x"9E9E9E9E",
		674 =>	x"9E9E9E9E",
		675 =>	x"9E9E9FA0",
		676 =>	x"9E9E9E9E",
		677 =>	x"9E9E9E9E",
		678 =>	x"9E9E9E9E",
		679 =>	x"9E9E9FA0",
		680 =>	x"9E9E9E9E",
		681 =>	x"9E9E9E9E",
		682 =>	x"9E9E9E9E",
		683 =>	x"9E9E9FA0",
		684 =>	x"9E9E9E9E",
		685 =>	x"9E9E9E9E",
		686 =>	x"9E9E9E9E",
		687 =>	x"9E9E9FA0",
		688 =>	x"9E9E9E9E",
		689 =>	x"9E9E9E9E",
		690 =>	x"9E9E9E9E",
		691 =>	x"9E9E9FA0",
		692 =>	x"9E9E9E9E",
		693 =>	x"9E9E9E9E",
		694 =>	x"9E9E9E9E",
		695 =>	x"9E9E9FA0",
		696 =>	x"9E9E9E9E",
		697 =>	x"9E9E9E9E",
		698 =>	x"9E9E9E9E",
		699 =>	x"9E9E9FA0",
		700 =>	x"9E9E9E9E",
		701 =>	x"9E9E9E9E",
		702 =>	x"9E9E9E9E",
		703 =>	x"9E9E9FA0",
		704 =>	x"A1A2A3A0", -- IMG_16x16_map_element_02
		705 =>	x"A0A0A0A0",
		706 =>	x"A0A0A0A0",
		707 =>	x"A0A0A0A0",
		708 =>	x"A4A5A6A7",
		709 =>	x"9F9F9F9F",
		710 =>	x"9F9F9F9F",
		711 =>	x"9F9F9F9F",
		712 =>	x"A3A89E9E",
		713 =>	x"9E9E9E9E",
		714 =>	x"9E9E9E9E",
		715 =>	x"9E9E9E9E",
		716 =>	x"A09F9E9E",
		717 =>	x"9E9E9E9E",
		718 =>	x"9E9E9E9E",
		719 =>	x"9E9E9E9E",
		720 =>	x"A09F9E9E",
		721 =>	x"9E9E9E9E",
		722 =>	x"9E9E9E9E",
		723 =>	x"9E9E9E9E",
		724 =>	x"A09F9E9E",
		725 =>	x"9E9E9E9E",
		726 =>	x"9E9E9E9E",
		727 =>	x"9E9E9E9E",
		728 =>	x"A09F9E9E",
		729 =>	x"9E9E9E9E",
		730 =>	x"9E9E9E9E",
		731 =>	x"9E9E9E9E",
		732 =>	x"A09F9E9E",
		733 =>	x"9E9E9E9E",
		734 =>	x"9E9E9E9E",
		735 =>	x"9E9E9E9E",
		736 =>	x"A09F9E9E",
		737 =>	x"9E9E9E9E",
		738 =>	x"9E9E9E9E",
		739 =>	x"9E9E9E9E",
		740 =>	x"A09F9E9E",
		741 =>	x"9E9E9E9E",
		742 =>	x"9E9E9E9E",
		743 =>	x"9E9E9E9E",
		744 =>	x"A09F9E9E",
		745 =>	x"9E9E9E9E",
		746 =>	x"9E9E9E9E",
		747 =>	x"9E9E9E9E",
		748 =>	x"A09F9E9E",
		749 =>	x"9E9E9E9E",
		750 =>	x"9E9E9E9E",
		751 =>	x"9E9E9E9E",
		752 =>	x"A09F9E9E",
		753 =>	x"9E9E9E9E",
		754 =>	x"9E9E9E9E",
		755 =>	x"9E9E9E9E",
		756 =>	x"A3A89E9E",
		757 =>	x"9E9E9E9E",
		758 =>	x"9E9E9E9E",
		759 =>	x"9E9E9E9E",
		760 =>	x"A4A5A6A7",
		761 =>	x"9F9F9F9F",
		762 =>	x"9F9F9F9F",
		763 =>	x"9F9F9F9F",
		764 =>	x"A1A2A3A0",
		765 =>	x"A0A0A0A0",
		766 =>	x"A0A0A0A0",
		767 =>	x"A0A0A0A0",
		768 =>	x"A09F9E9E", -- IMG_16x16_map_element_03
		769 =>	x"9E9E9E9E",
		770 =>	x"9E9E9E9E",
		771 =>	x"9E9E9FA0",
		772 =>	x"9FA99E9E",
		773 =>	x"9E9E9E9E",
		774 =>	x"9E9E9E9E",
		775 =>	x"9E9EA99F",
		776 =>	x"9E9E9E9E",
		777 =>	x"9E9E9E9E",
		778 =>	x"9E9E9E9E",
		779 =>	x"9E9E9E9E",
		780 =>	x"9E9E9E9E",
		781 =>	x"9E9E9E9E",
		782 =>	x"9E9E9E9E",
		783 =>	x"9E9E9E9E",
		784 =>	x"9E9E9E9E",
		785 =>	x"9E9E9E9E",
		786 =>	x"9E9E9E9E",
		787 =>	x"9E9E9E9E",
		788 =>	x"9E9E9E9E",
		789 =>	x"9E9E9E9E",
		790 =>	x"9E9E9E9E",
		791 =>	x"9E9E9E9E",
		792 =>	x"9E9E9E9E",
		793 =>	x"9E9E9E9E",
		794 =>	x"9E9E9E9E",
		795 =>	x"9E9E9E9E",
		796 =>	x"9E9E9E9E",
		797 =>	x"9E9E9E9E",
		798 =>	x"9E9E9E9E",
		799 =>	x"9E9E9E9E",
		800 =>	x"9E9E9E9E",
		801 =>	x"9E9E9E9E",
		802 =>	x"9E9E9E9E",
		803 =>	x"9E9E9E9E",
		804 =>	x"9E9E9E9E",
		805 =>	x"9E9E9E9E",
		806 =>	x"9E9E9E9E",
		807 =>	x"9E9E9E9E",
		808 =>	x"9E9E9E9E",
		809 =>	x"9E9E9E9E",
		810 =>	x"9E9E9E9E",
		811 =>	x"9E9E9E9E",
		812 =>	x"9E9E9E9E",
		813 =>	x"9E9E9E9E",
		814 =>	x"9E9E9E9E",
		815 =>	x"9E9E9E9E",
		816 =>	x"9E9E9E9E",
		817 =>	x"9E9E9E9E",
		818 =>	x"9E9E9E9E",
		819 =>	x"9E9E9E9E",
		820 =>	x"9E9E9E9E",
		821 =>	x"9E9E9E9E",
		822 =>	x"9E9E9E9E",
		823 =>	x"9E9E9E9E",
		824 =>	x"9FA99E9E",
		825 =>	x"9E9E9E9E",
		826 =>	x"9E9E9E9E",
		827 =>	x"9E9EA99F",
		828 =>	x"A09F9E9E",
		829 =>	x"9E9E9E9E",
		830 =>	x"9E9E9E9E",
		831 =>	x"9E9E9FA0",
		832 =>	x"A0A0A0A0", -- IMG_16x16_map_element_04
		833 =>	x"A0A0A0A0",
		834 =>	x"A0A0A0A0",
		835 =>	x"A0A3A2A1",
		836 =>	x"9F9F9F9F",
		837 =>	x"9F9F9F9F",
		838 =>	x"9F9F9F9F",
		839 =>	x"A7A6A5A4",
		840 =>	x"9E9E9E9E",
		841 =>	x"9E9E9E9E",
		842 =>	x"9E9E9E9E",
		843 =>	x"9E9EA8A3",
		844 =>	x"9E9E9E9E",
		845 =>	x"9E9E9E9E",
		846 =>	x"9E9E9E9E",
		847 =>	x"9E9E9FA0",
		848 =>	x"9E9E9E9E",
		849 =>	x"9E9E9E9E",
		850 =>	x"9E9E9E9E",
		851 =>	x"9E9E9FA0",
		852 =>	x"9E9E9E9E",
		853 =>	x"9E9E9E9E",
		854 =>	x"9E9E9E9E",
		855 =>	x"9E9E9FA0",
		856 =>	x"9E9E9E9E",
		857 =>	x"9E9E9E9E",
		858 =>	x"9E9E9E9E",
		859 =>	x"9E9E9FA0",
		860 =>	x"9E9E9E9E",
		861 =>	x"9E9E9E9E",
		862 =>	x"9E9E9E9E",
		863 =>	x"9E9E9FA0",
		864 =>	x"9E9E9E9E",
		865 =>	x"9E9E9E9E",
		866 =>	x"9E9E9E9E",
		867 =>	x"9E9E9FA0",
		868 =>	x"9E9E9E9E",
		869 =>	x"9E9E9E9E",
		870 =>	x"9E9E9E9E",
		871 =>	x"9E9E9FA0",
		872 =>	x"9E9E9E9E",
		873 =>	x"9E9E9E9E",
		874 =>	x"9E9E9E9E",
		875 =>	x"9E9E9FA0",
		876 =>	x"9E9E9E9E",
		877 =>	x"9E9E9E9E",
		878 =>	x"9E9E9E9E",
		879 =>	x"9E9E9FA0",
		880 =>	x"9E9E9E9E",
		881 =>	x"9E9E9E9E",
		882 =>	x"9E9E9E9E",
		883 =>	x"9E9E9FA0",
		884 =>	x"9E9E9E9E",
		885 =>	x"9E9E9E9E",
		886 =>	x"9E9E9E9E",
		887 =>	x"9E9EA8A3",
		888 =>	x"9F9F9F9F",
		889 =>	x"9F9F9F9F",
		890 =>	x"9F9F9F9F",
		891 =>	x"A7A6A5A4",
		892 =>	x"A0A0A0A0",
		893 =>	x"A0A0A0A0",
		894 =>	x"A0A0A0A0",
		895 =>	x"A0A3A2A1",
		896 =>	x"A09F9E9E", -- IMG_16x16_map_element_05
		897 =>	x"9E9E9E9E",
		898 =>	x"9E9E9E9E",
		899 =>	x"9E9E9E9E",
		900 =>	x"A09F9E9E",
		901 =>	x"9E9E9E9E",
		902 =>	x"9E9E9E9E",
		903 =>	x"9E9E9E9E",
		904 =>	x"A09F9E9E",
		905 =>	x"9E9E9E9E",
		906 =>	x"9E9E9E9E",
		907 =>	x"9E9E9E9E",
		908 =>	x"A09F9E9E",
		909 =>	x"9E9E9E9E",
		910 =>	x"9E9E9E9E",
		911 =>	x"9E9E9E9E",
		912 =>	x"A09F9E9E",
		913 =>	x"9E9E9E9E",
		914 =>	x"9E9E9E9E",
		915 =>	x"9E9E9E9E",
		916 =>	x"A09F9E9E",
		917 =>	x"9E9E9E9E",
		918 =>	x"9E9E9E9E",
		919 =>	x"9E9E9E9E",
		920 =>	x"A09F9E9E",
		921 =>	x"9E9E9E9E",
		922 =>	x"9E9E9E9E",
		923 =>	x"9E9E9E9E",
		924 =>	x"A09F9E9E",
		925 =>	x"9E9E9E9E",
		926 =>	x"9E9E9E9E",
		927 =>	x"9E9E9E9E",
		928 =>	x"A09F9E9E",
		929 =>	x"9E9E9E9E",
		930 =>	x"9E9E9E9E",
		931 =>	x"9E9E9E9E",
		932 =>	x"A09F9E9E",
		933 =>	x"9E9E9E9E",
		934 =>	x"9E9E9E9E",
		935 =>	x"9E9E9E9E",
		936 =>	x"A09F9E9E",
		937 =>	x"9E9E9E9E",
		938 =>	x"9E9E9E9E",
		939 =>	x"9E9E9E9E",
		940 =>	x"A09F9E9E",
		941 =>	x"9E9E9E9E",
		942 =>	x"9E9E9E9E",
		943 =>	x"9E9E9E9E",
		944 =>	x"A09F9E9E",
		945 =>	x"9E9E9E9E",
		946 =>	x"9E9E9E9E",
		947 =>	x"9E9E9E9E",
		948 =>	x"A3A89E9E",
		949 =>	x"9E9E9E9E",
		950 =>	x"9E9E9E9E",
		951 =>	x"9E9E9E9E",
		952 =>	x"A4A5A6A7",
		953 =>	x"9F9F9F9F",
		954 =>	x"9F9F9F9F",
		955 =>	x"9F9F9F9F",
		956 =>	x"A1A2A3A0",
		957 =>	x"A0A0A0A0",
		958 =>	x"A0A0A0A0",
		959 =>	x"A0A0A0A0",
		960 =>	x"9E9E9E9E", -- IMG_16x16_map_element_06
		961 =>	x"9E9E9E9E",
		962 =>	x"9E9E9E9E",
		963 =>	x"9E9E9E9E",
		964 =>	x"9E9E9E9E",
		965 =>	x"9E9E9E9E",
		966 =>	x"9E9E9E9E",
		967 =>	x"9E9E9E9E",
		968 =>	x"9E9E9E9E",
		969 =>	x"9E9E9E9E",
		970 =>	x"9E9E9E9E",
		971 =>	x"9E9E9E9E",
		972 =>	x"9E9E9E9E",
		973 =>	x"9E9E9E9E",
		974 =>	x"9E9E9E9E",
		975 =>	x"9E9E9E9E",
		976 =>	x"9E9E9E9E",
		977 =>	x"9E9E9E9E",
		978 =>	x"9E9E9E9E",
		979 =>	x"9E9E9E9E",
		980 =>	x"9E9E9E9E",
		981 =>	x"9E9E9E9E",
		982 =>	x"9E9E9E9E",
		983 =>	x"9E9E9E9E",
		984 =>	x"9E9E9E9E",
		985 =>	x"9E9E9E9E",
		986 =>	x"9E9E9E9E",
		987 =>	x"9E9E9E9E",
		988 =>	x"9E9E9E9E",
		989 =>	x"9E9E9E9E",
		990 =>	x"9E9E9E9E",
		991 =>	x"9E9E9E9E",
		992 =>	x"9E9E9E9E",
		993 =>	x"9E9E9E9E",
		994 =>	x"9E9E9E9E",
		995 =>	x"9E9E9E9E",
		996 =>	x"9E9E9E9E",
		997 =>	x"9E9E9E9E",
		998 =>	x"9E9E9E9E",
		999 =>	x"9E9E9E9E",
		1000 =>	x"9E9E9E9E",
		1001 =>	x"9E9E9E9E",
		1002 =>	x"9E9E9E9E",
		1003 =>	x"9E9E9E9E",
		1004 =>	x"9E9E9E9E",
		1005 =>	x"9E9E9E9E",
		1006 =>	x"9E9E9E9E",
		1007 =>	x"9E9E9E9E",
		1008 =>	x"9E9E9E9E",
		1009 =>	x"9E9E9E9E",
		1010 =>	x"9E9E9E9E",
		1011 =>	x"9E9E9E9E",
		1012 =>	x"9E9E9E9E",
		1013 =>	x"9E9E9E9E",
		1014 =>	x"9E9E9E9E",
		1015 =>	x"9E9E9E9E",
		1016 =>	x"9F9F9F9F",
		1017 =>	x"9F9F9F9F",
		1018 =>	x"9F9F9F9F",
		1019 =>	x"9F9F9F9F",
		1020 =>	x"A0A0A0A0",
		1021 =>	x"A0A0A0A0",
		1022 =>	x"A0A0A0A0",
		1023 =>	x"A0A0A0A0",
		1024 =>	x"9E9E9E9E", -- IMG_16x16_map_element_07
		1025 =>	x"9E9E9E9E",
		1026 =>	x"9E9E9E9E",
		1027 =>	x"9E9E9FA0",
		1028 =>	x"9E9E9E9E",
		1029 =>	x"9E9E9E9E",
		1030 =>	x"9E9E9E9E",
		1031 =>	x"9E9E9FA0",
		1032 =>	x"9E9E9E9E",
		1033 =>	x"9E9E9E9E",
		1034 =>	x"9E9E9E9E",
		1035 =>	x"9E9E9FA0",
		1036 =>	x"9E9E9E9E",
		1037 =>	x"9E9E9E9E",
		1038 =>	x"9E9E9E9E",
		1039 =>	x"9E9E9FA0",
		1040 =>	x"9E9E9E9E",
		1041 =>	x"9E9E9E9E",
		1042 =>	x"9E9E9E9E",
		1043 =>	x"9E9E9FA0",
		1044 =>	x"9E9E9E9E",
		1045 =>	x"9E9E9E9E",
		1046 =>	x"9E9E9E9E",
		1047 =>	x"9E9E9FA0",
		1048 =>	x"9E9E9E9E",
		1049 =>	x"9E9E9E9E",
		1050 =>	x"9E9E9E9E",
		1051 =>	x"9E9E9FA0",
		1052 =>	x"9E9E9E9E",
		1053 =>	x"9E9E9E9E",
		1054 =>	x"9E9E9E9E",
		1055 =>	x"9E9E9FA0",
		1056 =>	x"9E9E9E9E",
		1057 =>	x"9E9E9E9E",
		1058 =>	x"9E9E9E9E",
		1059 =>	x"9E9E9FA0",
		1060 =>	x"9E9E9E9E",
		1061 =>	x"9E9E9E9E",
		1062 =>	x"9E9E9E9E",
		1063 =>	x"9E9E9FA0",
		1064 =>	x"9E9E9E9E",
		1065 =>	x"9E9E9E9E",
		1066 =>	x"9E9E9E9E",
		1067 =>	x"9E9E9FA0",
		1068 =>	x"9E9E9E9E",
		1069 =>	x"9E9E9E9E",
		1070 =>	x"9E9E9E9E",
		1071 =>	x"9E9E9FA0",
		1072 =>	x"9E9E9E9E",
		1073 =>	x"9E9E9E9E",
		1074 =>	x"9E9E9E9E",
		1075 =>	x"9E9E9FA0",
		1076 =>	x"9E9E9E9E",
		1077 =>	x"9E9E9E9E",
		1078 =>	x"9E9E9E9E",
		1079 =>	x"9E9EA8A3",
		1080 =>	x"9F9F9F9F",
		1081 =>	x"9F9F9F9F",
		1082 =>	x"9F9F9F9F",
		1083 =>	x"A7A6A5A4",
		1084 =>	x"A0A0A0A0",
		1085 =>	x"A0A0A0A0",
		1086 =>	x"A0A0A0A0",
		1087 =>	x"A0A3A2A1",
		1088 =>	x"A09F9E9E", -- IMG_16x16_map_element_08
		1089 =>	x"9E9E9E9E",
		1090 =>	x"9E9E9E9E",
		1091 =>	x"9E9E9FA0",
		1092 =>	x"A09F9E9E",
		1093 =>	x"9E9E9E9E",
		1094 =>	x"9E9E9E9E",
		1095 =>	x"9E9EA99F",
		1096 =>	x"A09F9E9E",
		1097 =>	x"9E9E9E9E",
		1098 =>	x"9E9E9E9E",
		1099 =>	x"9E9E9E9E",
		1100 =>	x"A09F9E9E",
		1101 =>	x"9E9E9E9E",
		1102 =>	x"9E9E9E9E",
		1103 =>	x"9E9E9E9E",
		1104 =>	x"A09F9E9E",
		1105 =>	x"9E9E9E9E",
		1106 =>	x"9E9E9E9E",
		1107 =>	x"9E9E9E9E",
		1108 =>	x"A09F9E9E",
		1109 =>	x"9E9E9E9E",
		1110 =>	x"9E9E9E9E",
		1111 =>	x"9E9E9E9E",
		1112 =>	x"A09F9E9E",
		1113 =>	x"9E9E9E9E",
		1114 =>	x"9E9E9E9E",
		1115 =>	x"9E9E9E9E",
		1116 =>	x"A09F9E9E",
		1117 =>	x"9E9E9E9E",
		1118 =>	x"9E9E9E9E",
		1119 =>	x"9E9E9E9E",
		1120 =>	x"A09F9E9E",
		1121 =>	x"9E9E9E9E",
		1122 =>	x"9E9E9E9E",
		1123 =>	x"9E9E9E9E",
		1124 =>	x"A09F9E9E",
		1125 =>	x"9E9E9E9E",
		1126 =>	x"9E9E9E9E",
		1127 =>	x"9E9E9E9E",
		1128 =>	x"A09F9E9E",
		1129 =>	x"9E9E9E9E",
		1130 =>	x"9E9E9E9E",
		1131 =>	x"9E9E9E9E",
		1132 =>	x"A09F9E9E",
		1133 =>	x"9E9E9E9E",
		1134 =>	x"9E9E9E9E",
		1135 =>	x"9E9E9E9E",
		1136 =>	x"A09F9E9E",
		1137 =>	x"9E9E9E9E",
		1138 =>	x"9E9E9E9E",
		1139 =>	x"9E9E9E9E",
		1140 =>	x"A3A89E9E",
		1141 =>	x"9E9E9E9E",
		1142 =>	x"9E9E9E9E",
		1143 =>	x"9E9E9E9E",
		1144 =>	x"A4A5A6A7",
		1145 =>	x"9F9F9F9F",
		1146 =>	x"9F9F9F9F",
		1147 =>	x"9F9F9F9F",
		1148 =>	x"A1A2A3A0",
		1149 =>	x"A0A0A0A0",
		1150 =>	x"A0A0A0A0",
		1151 =>	x"A0A0A0A0",
		1152 =>	x"A09F9E9E", -- IMG_16x16_map_element_09
		1153 =>	x"9E9E9E9E",
		1154 =>	x"9E9E9E9E",
		1155 =>	x"9E9E9FA0",
		1156 =>	x"A09F9E9E",
		1157 =>	x"9E9E9E9E",
		1158 =>	x"9E9E9E9E",
		1159 =>	x"9E9E9FA0",
		1160 =>	x"A09F9E9E",
		1161 =>	x"9E9E9E9E",
		1162 =>	x"9E9E9E9E",
		1163 =>	x"9E9E9FA0",
		1164 =>	x"A09F9E9E",
		1165 =>	x"9E9E9E9E",
		1166 =>	x"9E9E9E9E",
		1167 =>	x"9E9E9FA0",
		1168 =>	x"A09F9E9E",
		1169 =>	x"9E9E9E9E",
		1170 =>	x"9E9E9E9E",
		1171 =>	x"9E9E9FA0",
		1172 =>	x"A09F9E9E",
		1173 =>	x"9E9E9E9E",
		1174 =>	x"9E9E9E9E",
		1175 =>	x"9E9E9FA0",
		1176 =>	x"A09F9E9E",
		1177 =>	x"9E9E9E9E",
		1178 =>	x"9E9E9E9E",
		1179 =>	x"9E9E9FA0",
		1180 =>	x"A09F9E9E",
		1181 =>	x"9E9E9E9E",
		1182 =>	x"9E9E9E9E",
		1183 =>	x"9E9E9FA0",
		1184 =>	x"A09F9E9E",
		1185 =>	x"9E9E9E9E",
		1186 =>	x"9E9E9E9E",
		1187 =>	x"9E9E9FA0",
		1188 =>	x"A09F9E9E",
		1189 =>	x"9E9E9E9E",
		1190 =>	x"9E9E9E9E",
		1191 =>	x"9E9E9FA0",
		1192 =>	x"A09F9E9E",
		1193 =>	x"9E9E9E9E",
		1194 =>	x"9E9E9E9E",
		1195 =>	x"9E9E9FA0",
		1196 =>	x"A09F9E9E",
		1197 =>	x"9E9E9E9E",
		1198 =>	x"9E9E9E9E",
		1199 =>	x"9E9E9FA0",
		1200 =>	x"A09F9E9E",
		1201 =>	x"9E9E9E9E",
		1202 =>	x"9E9E9E9E",
		1203 =>	x"9E9E9FA0",
		1204 =>	x"A3A89E9E",
		1205 =>	x"9E9E9E9E",
		1206 =>	x"9E9E9E9E",
		1207 =>	x"9E9EA8A3",
		1208 =>	x"A4A5A6A7",
		1209 =>	x"9F9F9F9F",
		1210 =>	x"9F9F9F9F",
		1211 =>	x"A7A6A5A4",
		1212 =>	x"A1A2A3A0",
		1213 =>	x"A0A0A0A0",
		1214 =>	x"A0A0A0A0",
		1215 =>	x"A0A3A2A1",
		1216 =>	x"A09F9E9E", -- IMG_16x16_map_element_10
		1217 =>	x"9E9E9E9E",
		1218 =>	x"9E9E9E9E",
		1219 =>	x"9E9E9FA0",
		1220 =>	x"9FA99E9E",
		1221 =>	x"9E9E9E9E",
		1222 =>	x"9E9E9E9E",
		1223 =>	x"9E9E9FA0",
		1224 =>	x"9E9E9E9E",
		1225 =>	x"9E9E9E9E",
		1226 =>	x"9E9E9E9E",
		1227 =>	x"9E9E9FA0",
		1228 =>	x"9E9E9E9E",
		1229 =>	x"9E9E9E9E",
		1230 =>	x"9E9E9E9E",
		1231 =>	x"9E9E9FA0",
		1232 =>	x"9E9E9E9E",
		1233 =>	x"9E9E9E9E",
		1234 =>	x"9E9E9E9E",
		1235 =>	x"9E9E9FA0",
		1236 =>	x"9E9E9E9E",
		1237 =>	x"9E9E9E9E",
		1238 =>	x"9E9E9E9E",
		1239 =>	x"9E9E9FA0",
		1240 =>	x"9E9E9E9E",
		1241 =>	x"9E9E9E9E",
		1242 =>	x"9E9E9E9E",
		1243 =>	x"9E9E9FA0",
		1244 =>	x"9E9E9E9E",
		1245 =>	x"9E9E9E9E",
		1246 =>	x"9E9E9E9E",
		1247 =>	x"9E9E9FA0",
		1248 =>	x"9E9E9E9E",
		1249 =>	x"9E9E9E9E",
		1250 =>	x"9E9E9E9E",
		1251 =>	x"9E9E9FA0",
		1252 =>	x"9E9E9E9E",
		1253 =>	x"9E9E9E9E",
		1254 =>	x"9E9E9E9E",
		1255 =>	x"9E9E9FA0",
		1256 =>	x"9E9E9E9E",
		1257 =>	x"9E9E9E9E",
		1258 =>	x"9E9E9E9E",
		1259 =>	x"9E9E9FA0",
		1260 =>	x"9E9E9E9E",
		1261 =>	x"9E9E9E9E",
		1262 =>	x"9E9E9E9E",
		1263 =>	x"9E9E9FA0",
		1264 =>	x"9E9E9E9E",
		1265 =>	x"9E9E9E9E",
		1266 =>	x"9E9E9E9E",
		1267 =>	x"9E9E9FA0",
		1268 =>	x"9E9E9E9E",
		1269 =>	x"9E9E9E9E",
		1270 =>	x"9E9E9E9E",
		1271 =>	x"9E9EA8A3",
		1272 =>	x"9F9F9F9F",
		1273 =>	x"9F9F9F9F",
		1274 =>	x"9F9F9F9F",
		1275 =>	x"A7A6A5A4",
		1276 =>	x"A0A0A0A0",
		1277 =>	x"A0A0A0A0",
		1278 =>	x"A0A0A0A0",
		1279 =>	x"A0A3A2A1",
		1280 =>	x"A1A2A3A0", -- IMG_16x16_map_element_11
		1281 =>	x"A0A0A0A0",
		1282 =>	x"A0A0A0A0",
		1283 =>	x"A0A0A0A0",
		1284 =>	x"A4A5A6A7",
		1285 =>	x"9F9F9F9F",
		1286 =>	x"9F9F9F9F",
		1287 =>	x"9F9F9F9F",
		1288 =>	x"A3A89E9E",
		1289 =>	x"9E9E9E9E",
		1290 =>	x"9E9E9E9E",
		1291 =>	x"9E9E9E9E",
		1292 =>	x"A09F9E9E",
		1293 =>	x"9E9E9E9E",
		1294 =>	x"9E9E9E9E",
		1295 =>	x"9E9E9E9E",
		1296 =>	x"A09F9E9E",
		1297 =>	x"9E9E9E9E",
		1298 =>	x"9E9E9E9E",
		1299 =>	x"9E9E9E9E",
		1300 =>	x"A09F9E9E",
		1301 =>	x"9E9E9E9E",
		1302 =>	x"9E9E9E9E",
		1303 =>	x"9E9E9E9E",
		1304 =>	x"A09F9E9E",
		1305 =>	x"9E9E9E9E",
		1306 =>	x"9E9E9E9E",
		1307 =>	x"9E9E9E9E",
		1308 =>	x"A09F9E9E",
		1309 =>	x"9E9E9E9E",
		1310 =>	x"9E9E9E9E",
		1311 =>	x"9E9E9E9E",
		1312 =>	x"A09F9E9E",
		1313 =>	x"9E9E9E9E",
		1314 =>	x"9E9E9E9E",
		1315 =>	x"9E9E9E9E",
		1316 =>	x"A09F9E9E",
		1317 =>	x"9E9E9E9E",
		1318 =>	x"9E9E9E9E",
		1319 =>	x"9E9E9E9E",
		1320 =>	x"A09F9E9E",
		1321 =>	x"9E9E9E9E",
		1322 =>	x"9E9E9E9E",
		1323 =>	x"9E9E9E9E",
		1324 =>	x"A09F9E9E",
		1325 =>	x"9E9E9E9E",
		1326 =>	x"9E9E9E9E",
		1327 =>	x"9E9E9E9E",
		1328 =>	x"A09F9E9E",
		1329 =>	x"9E9E9E9E",
		1330 =>	x"9E9E9E9E",
		1331 =>	x"9E9E9E9E",
		1332 =>	x"A09F9E9E",
		1333 =>	x"9E9E9E9E",
		1334 =>	x"9E9E9E9E",
		1335 =>	x"9E9E9E9E",
		1336 =>	x"A09F9E9E",
		1337 =>	x"9E9E9E9E",
		1338 =>	x"9E9E9E9E",
		1339 =>	x"9E9E9E9E",
		1340 =>	x"A09F9E9E",
		1341 =>	x"9E9E9E9E",
		1342 =>	x"9E9E9E9E",
		1343 =>	x"9E9E9E9E",
		1344 =>	x"A0A0A0A0", -- IMG_16x16_map_element_12
		1345 =>	x"A0A0A0A0",
		1346 =>	x"A0A0A0A0",
		1347 =>	x"A0A0A0A0",
		1348 =>	x"9F9F9F9F",
		1349 =>	x"9F9F9F9F",
		1350 =>	x"9F9F9F9F",
		1351 =>	x"9F9F9F9F",
		1352 =>	x"9E9E9E9E",
		1353 =>	x"9E9E9E9E",
		1354 =>	x"9E9E9E9E",
		1355 =>	x"9E9E9E9E",
		1356 =>	x"9E9E9E9E",
		1357 =>	x"9E9E9E9E",
		1358 =>	x"9E9E9E9E",
		1359 =>	x"9E9E9E9E",
		1360 =>	x"9E9E9E9E",
		1361 =>	x"9E9E9E9E",
		1362 =>	x"9E9E9E9E",
		1363 =>	x"9E9E9E9E",
		1364 =>	x"9E9E9E9E",
		1365 =>	x"9E9E9E9E",
		1366 =>	x"9E9E9E9E",
		1367 =>	x"9E9E9E9E",
		1368 =>	x"9E9E9E9E",
		1369 =>	x"9E9E9E9E",
		1370 =>	x"9E9E9E9E",
		1371 =>	x"9E9E9E9E",
		1372 =>	x"9E9E9E9E",
		1373 =>	x"9E9E9E9E",
		1374 =>	x"9E9E9E9E",
		1375 =>	x"9E9E9E9E",
		1376 =>	x"9E9E9E9E",
		1377 =>	x"9E9E9E9E",
		1378 =>	x"9E9E9E9E",
		1379 =>	x"9E9E9E9E",
		1380 =>	x"9E9E9E9E",
		1381 =>	x"9E9E9E9E",
		1382 =>	x"9E9E9E9E",
		1383 =>	x"9E9E9E9E",
		1384 =>	x"9E9E9E9E",
		1385 =>	x"9E9E9E9E",
		1386 =>	x"9E9E9E9E",
		1387 =>	x"9E9E9E9E",
		1388 =>	x"9E9E9E9E",
		1389 =>	x"9E9E9E9E",
		1390 =>	x"9E9E9E9E",
		1391 =>	x"9E9E9E9E",
		1392 =>	x"9E9E9E9E",
		1393 =>	x"9E9E9E9E",
		1394 =>	x"9E9E9E9E",
		1395 =>	x"9E9E9E9E",
		1396 =>	x"9E9E9E9E",
		1397 =>	x"9E9E9E9E",
		1398 =>	x"9E9E9E9E",
		1399 =>	x"9E9E9E9E",
		1400 =>	x"9FA99E9E",
		1401 =>	x"9E9E9E9E",
		1402 =>	x"9E9E9E9E",
		1403 =>	x"9E9EA99F",
		1404 =>	x"A09F9E9E",
		1405 =>	x"9E9E9E9E",
		1406 =>	x"9E9E9E9E",
		1407 =>	x"9E9E9FA0",
		1408 =>	x"A09F9E9E", -- IMG_16x16_map_element_13
		1409 =>	x"9E9E9E9E",
		1410 =>	x"9E9E9E9E",
		1411 =>	x"9E9E9FA0",
		1412 =>	x"A09F9E9E",
		1413 =>	x"9E9E9E9E",
		1414 =>	x"9E9E9E9E",
		1415 =>	x"9E9EA99F",
		1416 =>	x"A09F9E9E",
		1417 =>	x"9E9E9E9E",
		1418 =>	x"9E9E9E9E",
		1419 =>	x"9E9E9E9E",
		1420 =>	x"A09F9E9E",
		1421 =>	x"9E9E9E9E",
		1422 =>	x"9E9E9E9E",
		1423 =>	x"9E9E9E9E",
		1424 =>	x"A09F9E9E",
		1425 =>	x"9E9E9E9E",
		1426 =>	x"9E9E9E9E",
		1427 =>	x"9E9E9E9E",
		1428 =>	x"A09F9E9E",
		1429 =>	x"9E9E9E9E",
		1430 =>	x"9E9E9E9E",
		1431 =>	x"9E9E9E9E",
		1432 =>	x"A09F9E9E",
		1433 =>	x"9E9E9E9E",
		1434 =>	x"9E9E9E9E",
		1435 =>	x"9E9E9E9E",
		1436 =>	x"A09F9E9E",
		1437 =>	x"9E9E9E9E",
		1438 =>	x"9E9E9E9E",
		1439 =>	x"9E9E9E9E",
		1440 =>	x"A09F9E9E",
		1441 =>	x"9E9E9E9E",
		1442 =>	x"9E9E9E9E",
		1443 =>	x"9E9E9E9E",
		1444 =>	x"A09F9E9E",
		1445 =>	x"9E9E9E9E",
		1446 =>	x"9E9E9E9E",
		1447 =>	x"9E9E9E9E",
		1448 =>	x"A09F9E9E",
		1449 =>	x"9E9E9E9E",
		1450 =>	x"9E9E9E9E",
		1451 =>	x"9E9E9E9E",
		1452 =>	x"A09F9E9E",
		1453 =>	x"9E9E9E9E",
		1454 =>	x"9E9E9E9E",
		1455 =>	x"9E9E9E9E",
		1456 =>	x"A09F9E9E",
		1457 =>	x"9E9E9E9E",
		1458 =>	x"9E9E9E9E",
		1459 =>	x"9E9E9E9E",
		1460 =>	x"A09F9E9E",
		1461 =>	x"9E9E9E9E",
		1462 =>	x"9E9E9E9E",
		1463 =>	x"9E9E9E9E",
		1464 =>	x"A09F9E9E",
		1465 =>	x"9E9E9E9E",
		1466 =>	x"9E9E9E9E",
		1467 =>	x"9E9EA99F",
		1468 =>	x"A09F9E9E",
		1469 =>	x"9E9E9E9E",
		1470 =>	x"9E9E9E9E",
		1471 =>	x"9E9E9FA0",
		1472 =>	x"A09F9E9E", -- IMG_16x16_map_element_14
		1473 =>	x"9E9E9E9E",
		1474 =>	x"9E9E9E9E",
		1475 =>	x"9E9E9FA0",
		1476 =>	x"9FA99E9E",
		1477 =>	x"9E9E9E9E",
		1478 =>	x"9E9E9E9E",
		1479 =>	x"9E9EA99F",
		1480 =>	x"9E9E9E9E",
		1481 =>	x"9E9E9E9E",
		1482 =>	x"9E9E9E9E",
		1483 =>	x"9E9E9E9E",
		1484 =>	x"9E9E9E9E",
		1485 =>	x"9E9E9E9E",
		1486 =>	x"9E9E9E9E",
		1487 =>	x"9E9E9E9E",
		1488 =>	x"9E9E9E9E",
		1489 =>	x"9E9E9E9E",
		1490 =>	x"9E9E9E9E",
		1491 =>	x"9E9E9E9E",
		1492 =>	x"9E9E9E9E",
		1493 =>	x"9E9E9E9E",
		1494 =>	x"9E9E9E9E",
		1495 =>	x"9E9E9E9E",
		1496 =>	x"9E9E9E9E",
		1497 =>	x"9E9E9E9E",
		1498 =>	x"9E9E9E9E",
		1499 =>	x"9E9E9E9E",
		1500 =>	x"9E9E9E9E",
		1501 =>	x"9E9E9E9E",
		1502 =>	x"9E9E9E9E",
		1503 =>	x"9E9E9E9E",
		1504 =>	x"9E9E9E9E",
		1505 =>	x"9E9E9E9E",
		1506 =>	x"9E9E9E9E",
		1507 =>	x"9E9E9E9E",
		1508 =>	x"9E9E9E9E",
		1509 =>	x"9E9E9E9E",
		1510 =>	x"9E9E9E9E",
		1511 =>	x"9E9E9E9E",
		1512 =>	x"9E9E9E9E",
		1513 =>	x"9E9E9E9E",
		1514 =>	x"9E9E9E9E",
		1515 =>	x"9E9E9E9E",
		1516 =>	x"9E9E9E9E",
		1517 =>	x"9E9E9E9E",
		1518 =>	x"9E9E9E9E",
		1519 =>	x"9E9E9E9E",
		1520 =>	x"9E9E9E9E",
		1521 =>	x"9E9E9E9E",
		1522 =>	x"9E9E9E9E",
		1523 =>	x"9E9E9E9E",
		1524 =>	x"9E9E9E9E",
		1525 =>	x"9E9E9E9E",
		1526 =>	x"9E9E9E9E",
		1527 =>	x"9E9E9E9E",
		1528 =>	x"9F9F9F9F",
		1529 =>	x"9F9F9F9F",
		1530 =>	x"9F9F9F9F",
		1531 =>	x"9F9F9F9F",
		1532 =>	x"A0A0A0A0",
		1533 =>	x"A0A0A0A0",
		1534 =>	x"A0A0A0A0",
		1535 =>	x"A0A0A0A0",
		1536 =>	x"A09F9E9E", -- IMG_16x16_map_element_15
		1537 =>	x"9E9E9E9E",
		1538 =>	x"9E9E9E9E",
		1539 =>	x"9E9E9FA0",
		1540 =>	x"9FA99E9E",
		1541 =>	x"9E9E9E9E",
		1542 =>	x"9E9E9E9E",
		1543 =>	x"9E9E9FA0",
		1544 =>	x"9E9E9E9E",
		1545 =>	x"9E9E9E9E",
		1546 =>	x"9E9E9E9E",
		1547 =>	x"9E9E9FA0",
		1548 =>	x"9E9E9E9E",
		1549 =>	x"9E9E9E9E",
		1550 =>	x"9E9E9E9E",
		1551 =>	x"9E9E9FA0",
		1552 =>	x"9E9E9E9E",
		1553 =>	x"9E9E9E9E",
		1554 =>	x"9E9E9E9E",
		1555 =>	x"9E9E9FA0",
		1556 =>	x"9E9E9E9E",
		1557 =>	x"9E9E9E9E",
		1558 =>	x"9E9E9E9E",
		1559 =>	x"9E9E9FA0",
		1560 =>	x"9E9E9E9E",
		1561 =>	x"9E9E9E9E",
		1562 =>	x"9E9E9E9E",
		1563 =>	x"9E9E9FA0",
		1564 =>	x"9E9E9E9E",
		1565 =>	x"9E9E9E9E",
		1566 =>	x"9E9E9E9E",
		1567 =>	x"9E9E9FA0",
		1568 =>	x"9E9E9E9E",
		1569 =>	x"9E9E9E9E",
		1570 =>	x"9E9E9E9E",
		1571 =>	x"9E9E9FA0",
		1572 =>	x"9E9E9E9E",
		1573 =>	x"9E9E9E9E",
		1574 =>	x"9E9E9E9E",
		1575 =>	x"9E9E9FA0",
		1576 =>	x"9E9E9E9E",
		1577 =>	x"9E9E9E9E",
		1578 =>	x"9E9E9E9E",
		1579 =>	x"9E9E9FA0",
		1580 =>	x"9E9E9E9E",
		1581 =>	x"9E9E9E9E",
		1582 =>	x"9E9E9E9E",
		1583 =>	x"9E9E9FA0",
		1584 =>	x"9E9E9E9E",
		1585 =>	x"9E9E9E9E",
		1586 =>	x"9E9E9E9E",
		1587 =>	x"9E9E9FA0",
		1588 =>	x"9E9E9E9E",
		1589 =>	x"9E9E9E9E",
		1590 =>	x"9E9E9E9E",
		1591 =>	x"9E9E9FA0",
		1592 =>	x"9FA99E9E",
		1593 =>	x"9E9E9E9E",
		1594 =>	x"9E9E9E9E",
		1595 =>	x"9E9E9FA0",
		1596 =>	x"A09F9E9E",
		1597 =>	x"9E9E9E9E",
		1598 =>	x"9E9E9E9E",
		1599 =>	x"9E9E9FA0",
		1600 =>	x"A09F9E9E", -- IMG_16x16_map_element_16
		1601 =>	x"9E9E9E9E",
		1602 =>	x"9E9E9E9E",
		1603 =>	x"9E9E9FA0",
		1604 =>	x"A09F9E9E",
		1605 =>	x"9E9E9E9E",
		1606 =>	x"9E9E9E9E",
		1607 =>	x"9E9E9FA0",
		1608 =>	x"A09F9E9E",
		1609 =>	x"9E9E9E9E",
		1610 =>	x"9E9E9E9E",
		1611 =>	x"9E9E9FA0",
		1612 =>	x"A09F9E9E",
		1613 =>	x"9E9E9E9E",
		1614 =>	x"9E9E9E9E",
		1615 =>	x"9E9E9FA0",
		1616 =>	x"A09F9E9E",
		1617 =>	x"9E9E9E9E",
		1618 =>	x"9E9E9E9E",
		1619 =>	x"9E9E9FA0",
		1620 =>	x"A09F9E9E",
		1621 =>	x"9E9E9E9E",
		1622 =>	x"9E9E9E9E",
		1623 =>	x"9E9E9FA0",
		1624 =>	x"A09F9E9E",
		1625 =>	x"9E9E9E9E",
		1626 =>	x"9E9E9E9E",
		1627 =>	x"9E9E9FA0",
		1628 =>	x"A09F9E9E",
		1629 =>	x"9E9E9E9E",
		1630 =>	x"9E9E9E9E",
		1631 =>	x"9E9E9FA0",
		1632 =>	x"A09F9E9E",
		1633 =>	x"9E9E9E9E",
		1634 =>	x"9E9E9E9E",
		1635 =>	x"9E9E9FA0",
		1636 =>	x"A09F9E9E",
		1637 =>	x"9E9E9E9E",
		1638 =>	x"9E9E9E9E",
		1639 =>	x"9E9E9FA0",
		1640 =>	x"A09F9E9E",
		1641 =>	x"9E9E9E9E",
		1642 =>	x"9E9E9E9E",
		1643 =>	x"9E9E9FA0",
		1644 =>	x"A09F9E9E",
		1645 =>	x"9E9E9E9E",
		1646 =>	x"9E9E9E9E",
		1647 =>	x"9E9E9FA0",
		1648 =>	x"A09F9E9E",
		1649 =>	x"9E9E9E9E",
		1650 =>	x"9E9E9E9E",
		1651 =>	x"9E9E9FA0",
		1652 =>	x"A09F9E9E",
		1653 =>	x"9E9E9E9E",
		1654 =>	x"9E9E9E9E",
		1655 =>	x"9E9E9FA0",
		1656 =>	x"A09F9E9E",
		1657 =>	x"9E9E9E9E",
		1658 =>	x"9E9E9E9E",
		1659 =>	x"9E9E9FA0",
		1660 =>	x"A09F9E9E",
		1661 =>	x"9E9E9E9E",
		1662 =>	x"9E9E9E9E",
		1663 =>	x"9E9E9FA0",
		1664 =>	x"A0A0A0A0", -- IMG_16x16_map_element_17
		1665 =>	x"A0A0A0A0",
		1666 =>	x"A0A0A0A0",
		1667 =>	x"A0A0A0A0",
		1668 =>	x"9F9F9F9F",
		1669 =>	x"9F9F9F9F",
		1670 =>	x"9F9F9F9F",
		1671 =>	x"9F9F9F9F",
		1672 =>	x"9E9E9E9E",
		1673 =>	x"9E9E9E9E",
		1674 =>	x"9E9E9E9E",
		1675 =>	x"9E9E9E9E",
		1676 =>	x"9E9E9E9E",
		1677 =>	x"9E9E9E9E",
		1678 =>	x"9E9E9E9E",
		1679 =>	x"9E9E9E9E",
		1680 =>	x"9E9E9E9E",
		1681 =>	x"9E9E9E9E",
		1682 =>	x"9E9E9E9E",
		1683 =>	x"9E9E9E9E",
		1684 =>	x"9E9E9E9E",
		1685 =>	x"9E9E9E9E",
		1686 =>	x"9E9E9E9E",
		1687 =>	x"9E9E9E9E",
		1688 =>	x"9E9E9E9E",
		1689 =>	x"9E9E9E9E",
		1690 =>	x"9E9E9E9E",
		1691 =>	x"9E9E9E9E",
		1692 =>	x"9E9E9E9E",
		1693 =>	x"9E9E9E9E",
		1694 =>	x"9E9E9E9E",
		1695 =>	x"9E9E9E9E",
		1696 =>	x"9E9E9E9E",
		1697 =>	x"9E9E9E9E",
		1698 =>	x"9E9E9E9E",
		1699 =>	x"9E9E9E9E",
		1700 =>	x"9E9E9E9E",
		1701 =>	x"9E9E9E9E",
		1702 =>	x"9E9E9E9E",
		1703 =>	x"9E9E9E9E",
		1704 =>	x"9E9E9E9E",
		1705 =>	x"9E9E9E9E",
		1706 =>	x"9E9E9E9E",
		1707 =>	x"9E9E9E9E",
		1708 =>	x"9E9E9E9E",
		1709 =>	x"9E9E9E9E",
		1710 =>	x"9E9E9E9E",
		1711 =>	x"9E9E9E9E",
		1712 =>	x"9E9E9E9E",
		1713 =>	x"9E9E9E9E",
		1714 =>	x"9E9E9E9E",
		1715 =>	x"9E9E9E9E",
		1716 =>	x"9E9E9E9E",
		1717 =>	x"9E9E9E9E",
		1718 =>	x"9E9E9E9E",
		1719 =>	x"9E9E9E9E",
		1720 =>	x"9F9F9F9F",
		1721 =>	x"9F9F9F9F",
		1722 =>	x"9F9F9F9F",
		1723 =>	x"9F9F9F9F",
		1724 =>	x"A0A0A0A0",
		1725 =>	x"A0A0A0A0",
		1726 =>	x"A0A0A0A0",
		1727 =>	x"A0A0A0A0",
		1728 =>	x"A1A2A3A0", -- IMG_16x16_map_element_18
		1729 =>	x"A0A0A0A0",
		1730 =>	x"A0A0A0A0",
		1731 =>	x"A0A3A2A1",
		1732 =>	x"A4A5A6A7",
		1733 =>	x"9F9F9F9F",
		1734 =>	x"9F9F9F9F",
		1735 =>	x"9FAAABA2",
		1736 =>	x"A3A89E9E",
		1737 =>	x"9E9E9E9E",
		1738 =>	x"9E9E9E9E",
		1739 =>	x"9E9E9FA3",
		1740 =>	x"A09F9E9E",
		1741 =>	x"9E9E9E9E",
		1742 =>	x"9E9E9E9E",
		1743 =>	x"9E9E9FA0",
		1744 =>	x"A09F9E9E",
		1745 =>	x"9E9E9E9E",
		1746 =>	x"9E9E9E9E",
		1747 =>	x"9E9E9FA0",
		1748 =>	x"A09F9E9E",
		1749 =>	x"9E9E9E9E",
		1750 =>	x"9E9E9E9E",
		1751 =>	x"9E9E9FA0",
		1752 =>	x"A09F9E9E",
		1753 =>	x"9E9E9E9E",
		1754 =>	x"9E9E9E9E",
		1755 =>	x"9E9E9FA0",
		1756 =>	x"A09F9E9E",
		1757 =>	x"9E9E9E9E",
		1758 =>	x"9E9E9E9E",
		1759 =>	x"9E9E9FA0",
		1760 =>	x"A09F9E9E",
		1761 =>	x"9E9E9E9E",
		1762 =>	x"9E9E9E9E",
		1763 =>	x"9E9E9FA0",
		1764 =>	x"A09F9E9E",
		1765 =>	x"9E9E9E9E",
		1766 =>	x"9E9E9E9E",
		1767 =>	x"9E9E9FA0",
		1768 =>	x"A09F9E9E",
		1769 =>	x"9E9E9E9E",
		1770 =>	x"9E9E9E9E",
		1771 =>	x"9E9E9FA0",
		1772 =>	x"A09F9E9E",
		1773 =>	x"9E9E9E9E",
		1774 =>	x"9E9E9E9E",
		1775 =>	x"9E9E9FA0",
		1776 =>	x"A09F9E9E",
		1777 =>	x"9E9E9E9E",
		1778 =>	x"9E9E9E9E",
		1779 =>	x"9E9E9FA0",
		1780 =>	x"A39F9E9E",
		1781 =>	x"9E9E9E9E",
		1782 =>	x"9E9E9E9E",
		1783 =>	x"9E9E9FA3",
		1784 =>	x"A2ABAA9F",
		1785 =>	x"9F9F9F9F",
		1786 =>	x"9F9F9F9F",
		1787 =>	x"9FAAABA2",
		1788 =>	x"A1A2A3A0",
		1789 =>	x"A0A0A0A0",
		1790 =>	x"A0A0A0A0",
		1791 =>	x"A0A3A2A1",
		1792 =>	x"A0A0A0A0", -- IMG_16x16_map_element_19
		1793 =>	x"A0A0A0A0",
		1794 =>	x"A0A0A0A0",
		1795 =>	x"A0A0A0A0",
		1796 =>	x"9F9F9F9F",
		1797 =>	x"9F9F9F9F",
		1798 =>	x"9F9F9F9F",
		1799 =>	x"9F9F9F9F",
		1800 =>	x"9E9E9E9E",
		1801 =>	x"9E9E9E9E",
		1802 =>	x"9E9E9E9E",
		1803 =>	x"9E9E9E9E",
		1804 =>	x"9E9E9E9E",
		1805 =>	x"9E9E9E9E",
		1806 =>	x"9E9E9E9E",
		1807 =>	x"9E9E9E9E",
		1808 =>	x"9E9E9E9E",
		1809 =>	x"9E9E9E9E",
		1810 =>	x"9E9E9E9E",
		1811 =>	x"9E9E9E9E",
		1812 =>	x"9E9E9E9E",
		1813 =>	x"9E9E9E9E",
		1814 =>	x"9E9E9E9E",
		1815 =>	x"9E9E9E9E",
		1816 =>	x"9E9E9E9E",
		1817 =>	x"9E9E9E9E",
		1818 =>	x"9E9E9E9E",
		1819 =>	x"9E9E9E9E",
		1820 =>	x"9E9E9E9E",
		1821 =>	x"9E9E9E9E",
		1822 =>	x"9E9E9E9E",
		1823 =>	x"9E9E9E9E",
		1824 =>	x"9E9E9E9E",
		1825 =>	x"9E9E9E9E",
		1826 =>	x"9E9E9E9E",
		1827 =>	x"9E9E9E9E",
		1828 =>	x"9E9E9E9E",
		1829 =>	x"9E9E9E9E",
		1830 =>	x"9E9E9E9E",
		1831 =>	x"9E9E9E9E",
		1832 =>	x"9E9E9E9E",
		1833 =>	x"9E9E9E9E",
		1834 =>	x"9E9E9E9E",
		1835 =>	x"9E9E9E9E",
		1836 =>	x"9E9E9E9E",
		1837 =>	x"9E9E9E9E",
		1838 =>	x"9E9E9E9E",
		1839 =>	x"9E9E9E9E",
		1840 =>	x"9E9E9E9E",
		1841 =>	x"9E9E9E9E",
		1842 =>	x"9E9E9E9E",
		1843 =>	x"9E9E9E9E",
		1844 =>	x"9E9E9E9E",
		1845 =>	x"9E9E9E9E",
		1846 =>	x"9E9E9E9E",
		1847 =>	x"9E9E9E9E",
		1848 =>	x"9E9E9E9E",
		1849 =>	x"9E9E9E9E",
		1850 =>	x"9E9E9E9E",
		1851 =>	x"9E9E9E9E",
		1852 =>	x"9E9E9E9E",
		1853 =>	x"9E9E9E9E",
		1854 =>	x"9E9E9E9E",
		1855 =>	x"9E9E9E9E",
		1856 =>	x"A0A0A0A0", -- IMG_16x16_map_element_20
		1857 =>	x"A0A0A0A0",
		1858 =>	x"A0A0A0A0",
		1859 =>	x"A0A3A2A1",
		1860 =>	x"9F9F9F9F",
		1861 =>	x"9F9F9F9F",
		1862 =>	x"9F9F9F9F",
		1863 =>	x"A7A6A5A4",
		1864 =>	x"9E9E9E9E",
		1865 =>	x"9E9E9E9E",
		1866 =>	x"9E9E9E9E",
		1867 =>	x"9E9EA8A3",
		1868 =>	x"9E9E9E9E",
		1869 =>	x"9E9E9E9E",
		1870 =>	x"9E9E9E9E",
		1871 =>	x"9E9E9FA0",
		1872 =>	x"9E9E9E9E",
		1873 =>	x"9E9E9E9E",
		1874 =>	x"9E9E9E9E",
		1875 =>	x"9E9E9FA0",
		1876 =>	x"9E9E9E9E",
		1877 =>	x"9E9E9E9E",
		1878 =>	x"9E9E9E9E",
		1879 =>	x"9E9E9FA0",
		1880 =>	x"9E9E9E9E",
		1881 =>	x"9E9E9E9E",
		1882 =>	x"9E9E9E9E",
		1883 =>	x"9E9E9FA0",
		1884 =>	x"9E9E9E9E",
		1885 =>	x"9E9E9E9E",
		1886 =>	x"9E9E9E9E",
		1887 =>	x"9E9E9FA0",
		1888 =>	x"9E9E9E9E",
		1889 =>	x"9E9E9E9E",
		1890 =>	x"9E9E9E9E",
		1891 =>	x"9E9E9FA0",
		1892 =>	x"9E9E9E9E",
		1893 =>	x"9E9E9E9E",
		1894 =>	x"9E9E9E9E",
		1895 =>	x"9E9E9FA0",
		1896 =>	x"9E9E9E9E",
		1897 =>	x"9E9E9E9E",
		1898 =>	x"9E9E9E9E",
		1899 =>	x"9E9E9FA0",
		1900 =>	x"9E9E9E9E",
		1901 =>	x"9E9E9E9E",
		1902 =>	x"9E9E9E9E",
		1903 =>	x"9E9E9FA0",
		1904 =>	x"9E9E9E9E",
		1905 =>	x"9E9E9E9E",
		1906 =>	x"9E9E9E9E",
		1907 =>	x"9E9E9FA0",
		1908 =>	x"9E9E9E9E",
		1909 =>	x"9E9E9E9E",
		1910 =>	x"9E9E9E9E",
		1911 =>	x"9E9E9FA0",
		1912 =>	x"9E9E9E9E",
		1913 =>	x"9E9E9E9E",
		1914 =>	x"9E9E9E9E",
		1915 =>	x"9E9E9FA0",
		1916 =>	x"9E9E9E9E",
		1917 =>	x"9E9E9E9E",
		1918 =>	x"9E9E9E9E",
		1919 =>	x"9E9E9FA0",
		1920 =>	x"A1A2A3A0", -- IMG_16x16_map_element_21
		1921 =>	x"A0A0A0A0",
		1922 =>	x"A0A0A0A0",
		1923 =>	x"A0A0A0A0",
		1924 =>	x"A4A5A6A7",
		1925 =>	x"9F9F9F9F",
		1926 =>	x"9F9F9F9F",
		1927 =>	x"9F9F9F9F",
		1928 =>	x"A3A89E9E",
		1929 =>	x"9E9E9E9E",
		1930 =>	x"9E9E9E9E",
		1931 =>	x"9E9E9E9E",
		1932 =>	x"A09F9E9E",
		1933 =>	x"9E9E9E9E",
		1934 =>	x"9E9E9E9E",
		1935 =>	x"9E9E9E9E",
		1936 =>	x"A09F9E9E",
		1937 =>	x"9E9E9E9E",
		1938 =>	x"9E9E9E9E",
		1939 =>	x"9E9E9E9E",
		1940 =>	x"A09F9E9E",
		1941 =>	x"9E9E9E9E",
		1942 =>	x"9E9E9E9E",
		1943 =>	x"9E9E9E9E",
		1944 =>	x"A09F9E9E",
		1945 =>	x"9E9E9E9E",
		1946 =>	x"9E9E9E9E",
		1947 =>	x"9E9E9E9E",
		1948 =>	x"A09F9E9E",
		1949 =>	x"9E9E9E9E",
		1950 =>	x"9E9E9E9E",
		1951 =>	x"9E9E9E9E",
		1952 =>	x"A09F9E9E",
		1953 =>	x"9E9E9E9E",
		1954 =>	x"9E9E9E9E",
		1955 =>	x"9E9E9E9E",
		1956 =>	x"A09F9E9E",
		1957 =>	x"9E9E9E9E",
		1958 =>	x"9E9E9E9E",
		1959 =>	x"9E9E9E9E",
		1960 =>	x"A09F9E9E",
		1961 =>	x"9E9E9E9E",
		1962 =>	x"9E9E9E9E",
		1963 =>	x"9E9E9E9E",
		1964 =>	x"A09F9E9E",
		1965 =>	x"9E9E9E9E",
		1966 =>	x"9E9E9E9E",
		1967 =>	x"9E9E9E9E",
		1968 =>	x"A09F9E9E",
		1969 =>	x"9E9E9E9E",
		1970 =>	x"9E9E9E9E",
		1971 =>	x"9E9E9E9E",
		1972 =>	x"A09F9E9E",
		1973 =>	x"9E9E9E9E",
		1974 =>	x"9E9E9E9E",
		1975 =>	x"9E9E9E9E",
		1976 =>	x"A09F9E9E",
		1977 =>	x"9E9E9E9E",
		1978 =>	x"9E9E9E9E",
		1979 =>	x"9E9EA99F",
		1980 =>	x"A09F9E9E",
		1981 =>	x"9E9E9E9E",
		1982 =>	x"9E9E9E9E",
		1983 =>	x"9E9E9FA0",
		1984 =>	x"A1A2A3A0", -- IMG_16x16_map_element_22
		1985 =>	x"A0A0A0A0",
		1986 =>	x"A0A0A0A0",
		1987 =>	x"A0A3A2A1",
		1988 =>	x"A4A5A6A7",
		1989 =>	x"9F9F9F9F",
		1990 =>	x"9F9F9F9F",
		1991 =>	x"A7A6A5A4",
		1992 =>	x"A3A89E9E",
		1993 =>	x"9E9E9E9E",
		1994 =>	x"9E9E9E9E",
		1995 =>	x"9E9EA8A3",
		1996 =>	x"A09F9E9E",
		1997 =>	x"9E9E9E9E",
		1998 =>	x"9E9E9E9E",
		1999 =>	x"9E9E9FA0",
		2000 =>	x"A09F9E9E",
		2001 =>	x"9E9E9E9E",
		2002 =>	x"9E9E9E9E",
		2003 =>	x"9E9E9FA0",
		2004 =>	x"A09F9E9E",
		2005 =>	x"9E9E9E9E",
		2006 =>	x"9E9E9E9E",
		2007 =>	x"9E9E9FA0",
		2008 =>	x"A09F9E9E",
		2009 =>	x"9E9E9E9E",
		2010 =>	x"9E9E9E9E",
		2011 =>	x"9E9E9FA0",
		2012 =>	x"A09F9E9E",
		2013 =>	x"9E9E9E9E",
		2014 =>	x"9E9E9E9E",
		2015 =>	x"9E9E9FA0",
		2016 =>	x"A09F9E9E",
		2017 =>	x"9E9E9E9E",
		2018 =>	x"9E9E9E9E",
		2019 =>	x"9E9E9FA0",
		2020 =>	x"A09F9E9E",
		2021 =>	x"9E9E9E9E",
		2022 =>	x"9E9E9E9E",
		2023 =>	x"9E9E9FA0",
		2024 =>	x"A09F9E9E",
		2025 =>	x"9E9E9E9E",
		2026 =>	x"9E9E9E9E",
		2027 =>	x"9E9E9FA0",
		2028 =>	x"A09F9E9E",
		2029 =>	x"9E9E9E9E",
		2030 =>	x"9E9E9E9E",
		2031 =>	x"9E9E9FA0",
		2032 =>	x"A09F9E9E",
		2033 =>	x"9E9E9E9E",
		2034 =>	x"9E9E9E9E",
		2035 =>	x"9E9E9FA0",
		2036 =>	x"A09F9E9E",
		2037 =>	x"9E9E9E9E",
		2038 =>	x"9E9E9E9E",
		2039 =>	x"9E9E9FA0",
		2040 =>	x"A09F9E9E",
		2041 =>	x"9E9E9E9E",
		2042 =>	x"9E9E9E9E",
		2043 =>	x"9E9E9FA0",
		2044 =>	x"A09F9E9E",
		2045 =>	x"9E9E9E9E",
		2046 =>	x"9E9E9E9E",
		2047 =>	x"9E9E9FA0",
		2048 =>	x"A0A0A0A0", -- IMG_16x16_map_element_23
		2049 =>	x"A0A0A0A0",
		2050 =>	x"A0A0A0A0",
		2051 =>	x"A0A3A2A1",
		2052 =>	x"9F9F9F9F",
		2053 =>	x"9F9F9F9F",
		2054 =>	x"9F9F9F9F",
		2055 =>	x"A7A6A5A4",
		2056 =>	x"9E9E9E9E",
		2057 =>	x"9E9E9E9E",
		2058 =>	x"9E9E9E9E",
		2059 =>	x"9E9EA8A3",
		2060 =>	x"9E9E9E9E",
		2061 =>	x"9E9E9E9E",
		2062 =>	x"9E9E9E9E",
		2063 =>	x"9E9E9FA0",
		2064 =>	x"9E9E9E9E",
		2065 =>	x"9E9E9E9E",
		2066 =>	x"9E9E9E9E",
		2067 =>	x"9E9E9FA0",
		2068 =>	x"9E9E9E9E",
		2069 =>	x"9E9E9E9E",
		2070 =>	x"9E9E9E9E",
		2071 =>	x"9E9E9FA0",
		2072 =>	x"9E9E9E9E",
		2073 =>	x"9E9E9E9E",
		2074 =>	x"9E9E9E9E",
		2075 =>	x"9E9E9FA0",
		2076 =>	x"9E9E9E9E",
		2077 =>	x"9E9E9E9E",
		2078 =>	x"9E9E9E9E",
		2079 =>	x"9E9E9FA0",
		2080 =>	x"9E9E9E9E",
		2081 =>	x"9E9E9E9E",
		2082 =>	x"9E9E9E9E",
		2083 =>	x"9E9E9FA0",
		2084 =>	x"9E9E9E9E",
		2085 =>	x"9E9E9E9E",
		2086 =>	x"9E9E9E9E",
		2087 =>	x"9E9E9FA0",
		2088 =>	x"9E9E9E9E",
		2089 =>	x"9E9E9E9E",
		2090 =>	x"9E9E9E9E",
		2091 =>	x"9E9E9FA0",
		2092 =>	x"9E9E9E9E",
		2093 =>	x"9E9E9E9E",
		2094 =>	x"9E9E9E9E",
		2095 =>	x"9E9E9FA0",
		2096 =>	x"9E9E9E9E",
		2097 =>	x"9E9E9E9E",
		2098 =>	x"9E9E9E9E",
		2099 =>	x"9E9E9FA0",
		2100 =>	x"9E9E9E9E",
		2101 =>	x"9E9E9E9E",
		2102 =>	x"9E9E9E9E",
		2103 =>	x"9E9E9FA0",
		2104 =>	x"9FA99E9E",
		2105 =>	x"9E9E9E9E",
		2106 =>	x"9E9E9E9E",
		2107 =>	x"9E9E9FA0",
		2108 =>	x"A09F9E9E",
		2109 =>	x"9E9E9E9E",
		2110 =>	x"9E9E9E9E",
		2111 =>	x"9E9E9FA0",
		2112 =>	x"A09F9E9E", -- IMG_16x16_map_element_24
		2113 =>	x"9E9E9E9E",
		2114 =>	x"9E9E9E9E",
		2115 =>	x"9E9E9E9E",
		2116 =>	x"A09F9E9E",
		2117 =>	x"9E9E9E9E",
		2118 =>	x"9E9E9E9E",
		2119 =>	x"9E9E9E9E",
		2120 =>	x"A09F9E9E",
		2121 =>	x"9E9E9E9E",
		2122 =>	x"9E9E9E9E",
		2123 =>	x"9E9E9E9E",
		2124 =>	x"A09F9E9E",
		2125 =>	x"9E9E9E9E",
		2126 =>	x"9E9E9E9E",
		2127 =>	x"9E9E9E9E",
		2128 =>	x"A09F9E9E",
		2129 =>	x"9E9E9E9E",
		2130 =>	x"9E9E9E9E",
		2131 =>	x"9E9E9E9E",
		2132 =>	x"A09F9E9E",
		2133 =>	x"9E9E9E9E",
		2134 =>	x"9E9E9E9E",
		2135 =>	x"9E9E9E9E",
		2136 =>	x"A09F9E9E",
		2137 =>	x"9E9E9E9E",
		2138 =>	x"9E9E9E9E",
		2139 =>	x"9E9E9E9E",
		2140 =>	x"A09F9E9E",
		2141 =>	x"9E9E9E9E",
		2142 =>	x"9E9E9E9E",
		2143 =>	x"9E9E9E9E",
		2144 =>	x"A09F9E9E",
		2145 =>	x"9E9E9E9E",
		2146 =>	x"9E9E9E9E",
		2147 =>	x"9E9E9E9E",
		2148 =>	x"A09F9E9E",
		2149 =>	x"9E9E9E9E",
		2150 =>	x"9E9E9E9E",
		2151 =>	x"9E9E9E9E",
		2152 =>	x"A09F9E9E",
		2153 =>	x"9E9E9E9E",
		2154 =>	x"9E9E9E9E",
		2155 =>	x"9E9E9E9E",
		2156 =>	x"A09F9E9E",
		2157 =>	x"9E9E9E9E",
		2158 =>	x"9E9E9E9E",
		2159 =>	x"9E9E9E9E",
		2160 =>	x"A09F9E9E",
		2161 =>	x"9E9E9E9E",
		2162 =>	x"9E9E9E9E",
		2163 =>	x"9E9E9E9E",
		2164 =>	x"A09F9E9E",
		2165 =>	x"9E9E9E9E",
		2166 =>	x"9E9E9E9E",
		2167 =>	x"9E9E9E9E",
		2168 =>	x"A09F9E9E",
		2169 =>	x"9E9E9E9E",
		2170 =>	x"9E9E9E9E",
		2171 =>	x"9E9E9E9E",
		2172 =>	x"A09F9E9E",
		2173 =>	x"9E9E9E9E",
		2174 =>	x"9E9E9E9E",
		2175 =>	x"9E9E9E9E",
		2176 =>	x"9E9E9E9E", -- IMG_16x16_map_element_25
		2177 =>	x"9E9E9E9E",
		2178 =>	x"9E9E9E9E",
		2179 =>	x"9E9E9E9E",
		2180 =>	x"9E9E9E9E",
		2181 =>	x"9E9E9E9E",
		2182 =>	x"9E9E9E9E",
		2183 =>	x"9E9E9E9E",
		2184 =>	x"9E9E9E9E",
		2185 =>	x"9E9E9E9E",
		2186 =>	x"9E9E9E9E",
		2187 =>	x"9E9E9E9E",
		2188 =>	x"9E9E9E9E",
		2189 =>	x"9E9E9E9E",
		2190 =>	x"9E9E9E9E",
		2191 =>	x"9E9E9E9E",
		2192 =>	x"9E9E9E9E",
		2193 =>	x"9E9E9E9E",
		2194 =>	x"9E9E9E9E",
		2195 =>	x"9E9E9E9E",
		2196 =>	x"9E9E9E9E",
		2197 =>	x"9E9E9E9E",
		2198 =>	x"9E9E9E9E",
		2199 =>	x"9E9E9E9E",
		2200 =>	x"9E9E9E9E",
		2201 =>	x"9E9E9E9E",
		2202 =>	x"9E9E9E9E",
		2203 =>	x"9E9E9E9E",
		2204 =>	x"9E9E9E9E",
		2205 =>	x"9E9E9E9E",
		2206 =>	x"9E9E9E9E",
		2207 =>	x"9E9E9E9E",
		2208 =>	x"9E9E9E9E",
		2209 =>	x"9E9E9E9E",
		2210 =>	x"9E9E9E9E",
		2211 =>	x"9E9E9E9E",
		2212 =>	x"9E9E9E9E",
		2213 =>	x"9E9E9E9E",
		2214 =>	x"9E9E9E9E",
		2215 =>	x"9E9E9E9E",
		2216 =>	x"9E9E9E9E",
		2217 =>	x"9E9E9E9E",
		2218 =>	x"9E9E9E9E",
		2219 =>	x"9E9E9E9E",
		2220 =>	x"9E9E9E9E",
		2221 =>	x"9E9E9E9E",
		2222 =>	x"9E9E9E9E",
		2223 =>	x"9E9E9E9E",
		2224 =>	x"9E9E9E9E",
		2225 =>	x"9E9E9E9E",
		2226 =>	x"9E9E9E9E",
		2227 =>	x"9E9E9E9E",
		2228 =>	x"9E9E9E9E",
		2229 =>	x"9E9E9E9E",
		2230 =>	x"9E9E9E9E",
		2231 =>	x"9E9E9E9E",
		2232 =>	x"9E9E9E9E",
		2233 =>	x"9E9E9E9E",
		2234 =>	x"9E9E9E9E",
		2235 =>	x"9E9E9E9E",
		2236 =>	x"9E9E9E9E",
		2237 =>	x"9E9E9E9E",
		2238 =>	x"9E9E9E9E",
		2239 =>	x"9E9E9E9E",
		2240 =>	x"96969696", -- IMG_16x16_rock
		2241 =>	x"96969696",
		2242 =>	x"96969696",
		2243 =>	x"96969696",
		2244 =>	x"96969696",
		2245 =>	x"96000000",
		2246 =>	x"00009696",
		2247 =>	x"96969696",
		2248 =>	x"96969696",
		2249 =>	x"009B9B9B",
		2250 =>	x"9B9B0096",
		2251 =>	x"96969696",
		2252 =>	x"96969600",
		2253 =>	x"9B9B9B9B",
		2254 =>	x"9B9B0096",
		2255 =>	x"96969696",
		2256 =>	x"96960000",
		2257 =>	x"9B9B9B9B",
		2258 =>	x"9B000096",
		2259 =>	x"96969696",
		2260 =>	x"9696009B",
		2261 =>	x"9B000000",
		2262 =>	x"9B9B9B00",
		2263 =>	x"00000096",
		2264 =>	x"9600009B",
		2265 =>	x"9B9B9B00",
		2266 =>	x"9B9B9B9B",
		2267 =>	x"9B9B0000",
		2268 =>	x"009B0000",
		2269 =>	x"00009B00",
		2270 =>	x"9B9B9B00",
		2271 =>	x"9B9B9B00",
		2272 =>	x"009B9B9B",
		2273 =>	x"009B9B00",
		2274 =>	x"9B9B9B9B",
		2275 =>	x"009B0000",
		2276 =>	x"00009B9B",
		2277 =>	x"009B0000",
		2278 =>	x"9B009B9B",
		2279 =>	x"009B9B00",
		2280 =>	x"96009B9B",
		2281 =>	x"009B9B00",
		2282 =>	x"9B9B9B9B",
		2283 =>	x"9B9B0096",
		2284 =>	x"009B9B9B",
		2285 =>	x"009B9B9B",
		2286 =>	x"009B9B00",
		2287 =>	x"00000096",
		2288 =>	x"009B9B9B",
		2289 =>	x"9B9B9B00",
		2290 =>	x"009B0000",
		2291 =>	x"96969696",
		2292 =>	x"9600009B",
		2293 =>	x"9B9B9B00",
		2294 =>	x"9B9B9B00",
		2295 =>	x"96969696",
		2296 =>	x"9696009B",
		2297 =>	x"9B9B9B9B",
		2298 =>	x"9B9B0096",
		2299 =>	x"96969696",
		2300 =>	x"96969600",
		2301 =>	x"0000009B",
		2302 =>	x"00009696",
		2303 =>	x"96969696",
		2304 =>	x"96969696", -- IMG_16x16_smoke
		2305 =>	x"96969696",
		2306 =>	x"96969696",
		2307 =>	x"96969696",
		2308 =>	x"96969600",
		2309 =>	x"00000096",
		2310 =>	x"96969696",
		2311 =>	x"96000096",
		2312 =>	x"96960072",
		2313 =>	x"72720000",
		2314 =>	x"00000096",
		2315 =>	x"00727200",
		2316 =>	x"96007272",
		2317 =>	x"72720072",
		2318 =>	x"72727296",
		2319 =>	x"00727200",
		2320 =>	x"96000072",
		2321 =>	x"72727272",
		2322 =>	x"72727200",
		2323 =>	x"72727200",
		2324 =>	x"72727272",
		2325 =>	x"72000000",
		2326 =>	x"72720000",
		2327 =>	x"72720096",
		2328 =>	x"72727272",
		2329 =>	x"00727272",
		2330 =>	x"00727272",
		2331 =>	x"72727200",
		2332 =>	x"96727200",
		2333 =>	x"72727272",
		2334 =>	x"00000072",
		2335 =>	x"72727200",
		2336 =>	x"72727200",
		2337 =>	x"72727272",
		2338 =>	x"72720072",
		2339 =>	x"72727200",
		2340 =>	x"00727272",
		2341 =>	x"72727272",
		2342 =>	x"72720072",
		2343 =>	x"72729696",
		2344 =>	x"72727272",
		2345 =>	x"72727272",
		2346 =>	x"72720072",
		2347 =>	x"00000096",
		2348 =>	x"96007272",
		2349 =>	x"72727272",
		2350 =>	x"72720072",
		2351 =>	x"72727296",
		2352 =>	x"96007272",
		2353 =>	x"72727272",
		2354 =>	x"00727272",
		2355 =>	x"72720096",
		2356 =>	x"00727272",
		2357 =>	x"72007272",
		2358 =>	x"00727272",
		2359 =>	x"72720096",
		2360 =>	x"00000000",
		2361 =>	x"00007272",
		2362 =>	x"00727272",
		2363 =>	x"72000096",
		2364 =>	x"96969696",
		2365 =>	x"96960000",
		2366 =>	x"96960000",
		2367 =>	x"00969696",


--			***** MAP *****


		2368 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2369 =>	x"00000140", -- z: 0 rot: 0 ptr: 320
		2370 =>	x"00000180", -- z: 0 rot: 0 ptr: 384
		2371 =>	x"000001C0", -- z: 0 rot: 0 ptr: 448
		2372 =>	x"00000200", -- z: 0 rot: 0 ptr: 512
		2373 =>	x"00000240", -- z: 0 rot: 0 ptr: 576
		2374 =>	x"00000280", -- z: 0 rot: 0 ptr: 640
		2375 =>	x"000002C0", -- z: 0 rot: 0 ptr: 704
		2376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2377 =>	x"00000340", -- z: 0 rot: 0 ptr: 832
		2378 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2379 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2380 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2381 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2382 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2383 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2384 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2385 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2386 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2387 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2388 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2389 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2390 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2391 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2392 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2393 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2394 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2395 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2396 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2397 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2398 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2399 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2400 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2401 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2402 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2403 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2404 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2405 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2406 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2407 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2408 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2409 =>	x"00000380", -- z: 0 rot: 0 ptr: 896
		2410 =>	x"000003C0", -- z: 0 rot: 0 ptr: 960
		2411 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2412 =>	x"00000440", -- z: 0 rot: 0 ptr: 1088
		2413 =>	x"00000480", -- z: 0 rot: 0 ptr: 1152
		2414 =>	x"000004C0", -- z: 0 rot: 0 ptr: 1216
		2415 =>	x"00000500", -- z: 0 rot: 0 ptr: 1280
		2416 =>	x"00000540", -- z: 0 rot: 0 ptr: 1344
		2417 =>	x"00000580", -- z: 0 rot: 0 ptr: 1408
		2418 =>	x"000005C0", -- z: 0 rot: 0 ptr: 1472
		2419 =>	x"00000600", -- z: 0 rot: 0 ptr: 1536
		2420 =>	x"00000640", -- z: 0 rot: 0 ptr: 1600
		2421 =>	x"00000680", -- z: 0 rot: 0 ptr: 1664
		2422 =>	x"000006C0", -- z: 0 rot: 0 ptr: 1728
		2423 =>	x"00000700", -- z: 0 rot: 0 ptr: 1792
		2424 =>	x"00000740", -- z: 0 rot: 0 ptr: 1856
		2425 =>	x"000007C0", -- z: 0 rot: 0 ptr: 1984
		2426 =>	x"00000800", -- z: 0 rot: 0 ptr: 2048
		2427 =>	x"00000840", -- z: 0 rot: 0 ptr: 2112
		2428 =>	x"00000880", -- z: 0 rot: 0 ptr: 2176
		2429 =>	x"000004C0", -- z: 0 rot: 0 ptr: 1216
		2430 =>	x"00000600", -- z: 0 rot: 0 ptr: 1536
		2431 =>	x"000008C0", -- z: 0 rot: 0 ptr: 2240
		2432 =>	x"00000900", -- z: 0 rot: 0 ptr: 2304
		2433 =>	x"00000780", -- z: 0 rot: 0 ptr: 1920
		2434 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2435 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2436 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2437 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2438 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2439 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2440 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2441 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2442 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2443 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2444 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2445 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2446 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2447 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2448 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2449 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2450 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2451 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2452 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2453 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2454 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2455 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2456 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2457 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2458 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2459 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2460 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2461 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2462 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2463 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2464 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2465 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2466 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2467 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2468 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2469 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2470 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2471 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2472 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2473 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2474 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2475 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2476 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2477 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2478 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2479 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2480 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2481 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2482 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2483 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2484 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2485 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2486 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2487 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2488 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2489 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2490 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2491 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2492 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2493 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2494 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2495 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2496 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2497 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2498 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2499 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2500 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2501 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2502 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2503 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2504 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2505 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2506 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2507 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2508 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2509 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2510 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2511 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2512 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2513 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2514 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2515 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2516 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2517 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2518 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2519 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2520 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2521 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2522 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2523 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2524 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2525 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2526 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2527 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2528 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2529 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2530 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2531 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2532 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2533 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2534 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2535 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2536 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2537 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2538 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2539 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2540 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2541 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2542 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2543 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2544 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2545 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2546 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2547 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2548 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2549 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2550 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2551 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2552 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2553 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2554 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2555 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2556 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2557 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2558 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2559 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2560 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2561 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2562 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2563 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2564 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2565 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2566 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2567 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2568 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2569 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2570 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2571 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2572 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2573 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2574 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2575 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2576 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2577 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2578 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2579 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2580 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2581 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2582 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2583 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2584 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2585 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2586 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2587 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2588 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2589 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2590 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2591 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2592 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2593 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2594 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2595 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2596 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2597 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2598 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2599 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2600 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2601 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2602 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2603 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2604 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2605 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2606 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2607 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2608 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2609 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2610 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2611 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2612 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2613 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2614 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2615 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2616 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2617 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2618 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2619 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2620 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2621 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2622 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2623 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2624 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2625 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2626 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2627 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2628 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2629 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2630 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2631 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2632 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2633 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2634 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2635 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2636 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2637 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2638 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2639 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2640 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2641 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2642 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2643 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2644 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2645 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2646 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2647 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2648 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2649 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2650 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2651 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2652 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2653 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2654 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2655 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2656 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2657 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2658 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2659 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2660 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2661 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2662 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2663 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2664 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2665 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2666 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2667 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2668 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2669 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2670 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2671 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2672 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2673 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2674 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2675 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2676 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2677 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2678 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2679 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2680 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2681 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2682 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2683 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2684 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2685 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2686 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2687 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2688 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2689 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2690 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2691 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2692 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2693 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2694 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2695 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2696 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2697 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2698 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2699 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2700 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2701 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2702 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2703 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2704 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2705 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2706 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2707 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2708 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2709 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2710 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2711 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2712 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2713 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2714 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2715 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2716 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2717 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2718 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2719 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2720 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2721 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2722 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2723 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2724 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2725 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2726 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2727 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2728 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2729 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2730 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2731 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2732 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2733 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2734 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2735 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2736 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2737 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2738 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2739 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2740 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2741 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2742 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2743 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2744 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2745 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2746 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2747 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2748 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2749 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2750 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2751 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2752 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2753 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2754 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2755 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2756 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2757 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2758 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2759 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2760 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2761 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2762 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2763 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2764 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2765 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2766 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2767 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2768 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2769 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2770 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2771 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2772 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2773 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2774 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2775 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2776 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2777 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2778 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2779 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2780 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2781 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2782 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2783 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2784 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2785 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2786 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2787 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2788 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2789 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2790 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2791 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2792 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2793 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2794 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2795 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2796 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2797 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2798 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2799 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2800 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2801 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2802 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2803 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2804 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2805 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2806 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2807 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2808 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2809 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2810 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2811 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2812 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2813 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2814 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2815 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2816 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2817 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2818 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2819 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2820 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2821 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2822 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2823 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2824 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2825 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2826 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2827 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2828 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2829 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2830 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2831 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2832 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2833 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2834 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2835 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2836 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2837 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2838 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2839 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2840 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2841 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2842 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2843 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2844 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2845 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2846 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2847 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2848 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2849 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2850 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2851 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2852 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2853 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2854 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2855 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2856 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2857 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2858 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2859 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2860 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2861 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2862 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2863 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2864 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2865 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2866 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2867 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2868 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2869 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2870 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2871 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2872 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2873 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2874 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2875 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2876 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2877 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2878 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2879 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2880 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2881 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2882 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2883 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2884 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2885 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2886 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2887 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2888 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2889 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2890 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2891 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2892 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2893 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2894 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2895 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2896 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2897 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2898 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2899 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2900 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2901 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2902 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2903 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2904 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2905 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2906 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2907 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2908 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2909 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2910 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2911 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2912 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2913 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2914 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2915 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2916 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2917 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2918 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2919 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2920 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2921 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2922 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2923 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2924 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2925 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2926 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2927 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2928 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2929 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2930 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2931 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2932 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2933 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2934 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2935 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2936 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2937 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2938 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2939 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2940 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2941 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2942 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2943 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2944 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2945 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2946 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2947 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2948 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2949 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2950 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2951 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2952 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2953 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2954 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2955 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2956 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2957 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2958 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2959 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2960 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2961 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2962 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2963 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2964 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2965 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2966 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2967 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2968 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2969 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2970 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2971 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2972 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2973 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2974 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2975 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2976 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2977 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2978 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2979 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2980 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2981 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2982 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2983 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2984 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2985 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2986 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2987 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2988 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2989 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2990 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2991 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2992 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2993 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2994 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2995 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2996 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2997 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2998 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2999 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3000 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3001 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3002 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3003 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3004 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3005 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3006 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3007 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3008 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3009 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3010 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3011 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3012 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3013 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3014 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3015 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3016 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3017 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3018 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3019 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3020 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3021 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3022 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3023 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3024 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3025 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3026 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3027 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3028 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3029 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3030 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3031 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3032 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3033 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3034 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3035 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3036 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3037 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3038 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3039 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3040 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3041 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3042 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3043 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3044 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3045 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3046 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3047 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3048 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3049 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3050 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3051 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3052 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3053 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3054 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3055 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3056 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3057 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3058 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3059 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3060 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3061 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3062 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3063 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3064 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3065 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3066 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3067 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3068 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3069 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3070 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3071 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3072 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3073 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3074 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3075 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3076 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3077 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3078 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3079 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3080 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3081 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3082 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3083 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3084 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3085 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3086 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3087 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3088 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3089 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3090 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3091 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3092 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3093 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3094 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3095 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3096 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3097 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3098 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3099 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3100 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3101 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3102 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3103 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3104 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3105 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3106 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3107 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3108 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3109 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3110 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3111 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3112 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3113 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3114 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3115 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3116 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3117 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3118 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3119 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3120 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3121 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3122 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3123 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3124 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3125 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3126 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3127 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3128 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3129 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3130 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3131 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3132 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3133 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3134 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3135 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3136 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3137 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3138 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3139 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3140 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3141 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3142 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3143 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3144 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3145 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3146 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3147 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3148 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3149 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3150 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3151 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3152 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3153 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3154 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3155 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3156 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3157 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3158 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3159 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3160 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3161 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3162 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3163 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3164 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3165 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3166 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3167 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3168 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3169 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3170 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3171 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3172 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3173 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3174 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3175 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3176 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3177 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3178 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3179 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3180 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3181 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3182 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3183 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3184 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3185 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3186 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3187 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3188 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3189 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3190 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3191 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3192 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3193 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3194 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3195 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3196 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3197 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3198 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3199 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3200 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3201 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3202 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3203 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3204 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3205 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3206 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3207 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3208 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3209 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3210 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3211 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3212 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3213 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3214 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3215 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3216 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3217 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3218 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3219 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3220 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3221 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3222 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3223 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3224 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3225 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3226 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3227 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3228 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3229 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3230 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3231 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3232 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3233 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3234 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3235 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3236 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3237 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3238 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3239 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3240 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3241 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3242 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3243 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3244 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3245 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3246 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3247 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3248 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3249 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3250 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3251 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3252 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3253 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3254 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3255 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3256 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3257 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3258 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3259 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3260 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3261 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3262 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3263 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3264 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3265 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3266 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3267 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3268 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3269 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3270 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3271 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3272 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3273 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3274 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3275 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3276 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3277 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3278 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3279 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3280 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3281 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3282 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3283 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3284 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3285 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3286 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3287 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3288 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3289 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3290 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3291 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3292 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3293 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3294 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3295 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3296 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3297 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3298 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3299 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3300 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3301 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3302 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3303 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3304 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3305 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3306 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3307 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3308 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3309 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3310 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3311 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3312 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3313 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3314 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3315 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3316 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3317 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3318 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3319 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3320 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3321 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3322 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3323 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3324 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3325 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3326 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3327 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3328 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3329 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3330 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3331 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3332 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3333 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3334 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3335 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3336 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3337 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3338 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3339 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3340 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3341 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3342 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3343 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3344 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3345 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3346 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3347 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3348 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3349 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3350 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3351 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3352 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3353 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3354 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3355 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3356 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3357 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3358 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3359 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3360 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3361 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3362 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3363 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3364 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3365 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3366 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3367 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3368 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3369 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3370 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3371 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3372 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3373 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3374 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3375 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3376 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3377 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3378 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3379 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3380 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3381 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3382 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3383 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3384 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3385 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3386 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3387 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3388 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3389 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3390 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3391 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3392 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3393 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3394 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3395 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3396 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3397 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3398 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3399 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3400 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3401 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3402 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3403 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3404 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3405 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3406 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3407 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3408 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3409 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3410 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3411 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3412 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3413 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3414 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3415 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3416 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3417 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3418 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3419 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3420 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3421 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3422 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3423 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3424 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3425 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3426 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3427 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3428 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3429 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3430 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3431 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3432 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3433 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3434 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3435 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3436 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3437 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3438 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3439 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3440 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3441 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3442 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3443 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3444 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3445 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3446 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3447 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3448 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3449 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3450 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3451 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3452 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3453 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3454 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3455 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3456 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3457 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3458 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3459 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3460 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3461 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3462 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3463 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3464 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3465 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3466 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3467 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3468 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3469 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3470 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3471 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3472 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3473 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3474 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3475 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3476 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3477 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3478 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3479 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3480 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3481 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3482 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3483 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3484 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3485 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3486 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3487 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3488 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3489 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3490 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3491 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3492 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3493 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3494 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3495 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3496 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3497 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3498 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3499 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3500 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3501 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3502 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3503 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3504 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3505 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3506 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3507 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3508 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3509 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3510 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3511 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3512 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3513 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3514 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3515 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3516 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3517 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3518 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3519 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3520 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3521 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3522 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3523 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3524 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3525 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3526 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3527 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3528 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3529 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3530 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3531 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3532 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3533 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3534 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3535 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3536 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3537 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3538 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3539 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3540 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3541 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3542 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3543 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3544 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3545 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3546 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3547 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3548 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3549 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3550 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3551 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3552 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3553 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3554 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3555 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3556 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3557 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3558 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3559 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3560 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3561 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3562 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3563 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3564 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3565 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3566 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3567 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3568 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3569 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3570 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3571 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3572 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3573 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3574 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3575 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3576 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3577 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3578 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3579 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3580 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3581 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3582 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3583 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3584 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3585 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3586 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3587 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3588 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3589 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3590 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3591 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3592 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3593 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3594 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3595 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3596 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3597 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3598 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3599 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3600 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3601 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3602 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3603 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3604 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3605 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3606 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3607 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3608 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3609 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3610 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3611 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3612 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3613 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3614 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3615 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3616 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3617 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3618 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3619 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3620 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3621 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3622 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3623 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3624 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3625 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3626 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3627 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3628 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3629 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3630 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3631 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3632 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3633 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3634 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3635 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3636 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3637 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3638 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		others => x"00000000"
	);

begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;